-- (C) 2001-2016 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
1twCu44N6z+K4X0ytMZzw/RrBml5HcQq69GDocLeINWP6oqYzwRUcKTFfIq/TCrkhPHCnnQ03Bgg
sx86Btti2C8lYfLAkQ5QjzN44VTqDFQaYY7DF0cvDNdcFnF9ZX0wyDU/gGggP/VzVuH4qA4ZvyHH
Puj/XJvQCWte00zh6k7DXGYuZPHFbWv1I67QxwHtoq6DyymfwHNW3LQWnER1QlvTKb2pOG6wOfMN
BpDIIHMMtCbfZKp4zpz2I+SqAhLM10zRN1NJSpr71i9FIqMTSHDTGxFjbLfP6Iokn2vlBnl6/cyG
SWXYmu4gyFgGf/mXDxY6HI9Ial8OQ2Uyb2ZeQQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 17344)
`protect data_block
CNqvih96WnkMORAY/U45BdlrjBZ8zKqCSJqwAqQI4CcVIcXTSTGB/vuqBMpmPues7owd0CIvVisz
8lX8GRU6GEyLwAjc9GO921/c8r8ITf7mP9VSH/nSlBpShUaDRfo+tP/+ukN6e85WjqnAuTL8cpoi
cQz2gDt+xL2CKtUGoWRr7DpoUh0fKAdIs0rbhf85U7Pf9ry27vz+yksXBwjk0sK3ieojQb2vJ4af
TrvDD9R7DyF4R/MKH78KjuDzwEJG+VwDHsf3fmJM+AuScXYsADDMf8oQhErEaNm2ee5nAfBKhGCm
WELrm3Yz0BtOKASpatZy2U8oHGtOZI7VZN9XaMWZuXxFaX+p07SSTq/fdxaV+1igJ21b5CvtujBc
qId8MloXErsxOpw7zEyIfoU3yOVUKZG3hCgxycAoyBv249ebot9JzP6y3Gp6Gbl/I1ELo13dIyUQ
jt3FedzJeP/WeyHfsm7ztJnZlZKVXeDioCJQ75WiblhDa5wPV7ZeNgrNWkDcSEfCaMgSUzMFu48v
Dkc2S/ydGVfVWLIAsUMHutw7HNkbTk9PHU9ptWymXdyzQXhYA49AmvwrkyojQpukEgzKngbsz80B
H7gw1Zv/24YGD2CxmZnDns65aqt6YZJSch4ZKBSxPtK5XxA2dWIAVNHQ/U/jBs36xQMnTQ339vAV
D0KPinBT5aBi5n2yAauPUuzcPJy0ckLMVUGNy4nLNaIkzy7adn72zipeLPk+fEw1obAxR+9myVYd
jn85q3CN/FZLcvONaIZk58eOFOHu6tYX69S0d1grYhqix3+NTW5+5DoKhbOxptPR/Thu7m9XllI2
fGEePxiCEDIjF279JI92einIP3we7XkMenFcuCM7YngWwuZniSSa7UvoEuGt5prDAYCeh8fGv8fT
XjReQpCSvWrMU1QfzsWwdRJGO/G+xxj+Ug34MoA65WHn6z+zwMiUwm4XtJ+WQ/skkQUZ9IpdX6dx
NNxCrazH/RUpp5id6N5mfcU/QrxH2EEpeVxw+SVkIY17ONnw0+WUfyL0+7wwiQ+r8MWtkfY4OAZY
W17LsIFGY25rgMMp0VMiY2X/pm6kl8JYb/m991n1PaGzy9vECvzEYf3X0TENXxTX1p9U5GFITAEL
hkesnPeSeNkKNmpym/Dn4vzw8VogTi8gHtGsGHaUPgg0oc02nCWtV88shHIrR1mcsNHfurPVVZbi
s7pvPiEwGFJOVB3hga9DobIho5kc3B7+zgMIBKX9N1xC/B/71zJ+saoWml9CsPIYg3G2yA4s15OO
mp3wBtKAQg3RI+1692BcIbelWqVOQwlwHcjX1dpnh6DROsUHaJK7RJKA87SZVsUAB4fIyW3fxLq7
MzVktxLPeONXqSiCCqFQVNUFQDsBP569FVzTaHE0/9fq2dMOt9PSDp2opb7vQoC6t7VwUVYhWLe3
EuJtzSbu3Y59AzE24TMdlVPn0Wq2bJBsb99Q82ndg3tiuJo1vIuqylJFePwU/DqwQi+l8gJr0IF2
IESz0TFrmQyIGFmHnOipjfNgcRH7UuuKaF5eDf6CvNBwcaxcfqsW8VgpqPLg75FLhIJegRMhRd1g
1OtDH1bz+CNJbE0ZK4ETEplgV2tbtL7ZFS8g2cCdCyXIySadqygn2idQzf0aIlx4ZGKpKhMfAEca
6A+iHiiK1unU8kUUBiCtpuFM3r4sZ5Q45O0Ljnfddt8CNwmzxmIFnnx5bZ8dt/Q9fyrQwYrcY2GH
7/9lc1fjMOFHMIiFoksWLUGLNIMP4kYVQXo7380dYyX3mfsqqgo0cnZa33WTmw3oJ9AaiT3JlohW
npOJT12YK/FO/j3pajhB7p80qsMH1mUJyCs1tgDHCR3fVkQ4dNmIdmhP+H/GrL5l5xV1OxTeA41Y
cWJg9UG2Ptva2PNzkAOfQnlFWUKHEkPutsOxWMhi6FG+8pYYQwYx9FmOR6UOyxbUZjRjudT62Mg/
eON7qIYFFSdjCqJuQKRYEXhoaF2OHtl0xAARTFk81n7sjTdJzKqZyG6IrH+st7+tsBvfGB97UsSD
zBZ9yk/5qRMPJ3sMiLHCUwE23+R9SYShLwq2jLHS1YrlOGVLV/h4kVfBMsk+g1Bmlni/7Vsu0Fqy
ZO+mVZVoWJEYpAltR4mykP1iDKm/JpunH1umdLShk5s/fiAm5O+l/VdPr2mT9T/tm2aWEvPpTNg6
VmIYJCLA17pCBKU3s7jRVU13+KiG+qZPCpBYfcpGgzCcXqG43ZKkO/nT7UmWR1EjQfyN+RouhNMx
q2hO33qEr7uaLEeqpKf/acFiQPdinuwfX1ggrzO78L3tQtoKQifQz5WT2ZFh+ZufO7Jyzf3biV+1
epsBGsfEoAFfcmF8X6QKV48VJGYDo5cBjJ6zHxEJX8NRULMVSMWu3otrqxYz1/S4f4R9Kwoh7Bse
28FbsLVErZ3KxRD16HASNt1wjNTvE4S5doHGo1IkEJUA9sb+XTMTaHG0kl1ur/BlDTdB0I9h5up/
lRIRhaxTNdz1IocjSQV8narc9BYLnjFeHSCVSqd89kUZoTQRuLmyqv3UwH21FWpD+D7lJJ4LJjUr
ia3VCc/F6VO32uHUdmPqBIowBb37rkhfyonmlXv7GwQPcQomytpFUo44Z7bDyVX2gkD1ohSycAEQ
v5ka60/T3e5maJ4Ck27R7vxLYgyj+ZmaQu+z7Elke49yBxk1APCMk21A2NQKrTggAkGaUHt8jHjR
UYXENeH8w7zQkDhJBhItP/1y+LIdQEEdGWww8cJJfWgHIBYIUnHmQINLjMsPdXMxSD5Q2g7Y2IYE
OUvmDoi7CBR0A71O3XyE2t8OPVbi3xyy4rOOnsmreYZp2KLP9w/2SKNQ1SjMPQzsh92uHx1fONJ8
GwTaRkO0gchQ6/8b6wN/h7wEpgNtkEYbuxzPR3V1sXq6oNsyMpRZSgZ9bWRWJ1xZowo+xD+4GX7F
YZgZgjT1HQmgAlQbiW40NrAGOlqzThiqJaaKnQ0BWWpHur/VfivxDTMbekzOcZc//tLO4QrbPg/n
sH+MkK6ImU8zFMKxgzN4uyY1DGhV/V9jG5dMyBhxdcz9Y69qOVQG8sUe3b59Kpb1E6A92cvkDqP+
xWOFu1WEDpwG0xOiNE/qzbFM1h54pOnw3dMvQ8l/IOhm2kktZ17Al+dCaX4BJO8t+9BaxJPKBE34
Coe1qBPvFbGTez+O9vWUomllLub9tbBcYjyiVTPqsLS1sboW/TTUcn08mxDb9Av2u+6O4wBsKa14
UoVo5+IgKevdnw7RiS/HGCEifNDko4PL9YcpfoEh36in9oHY/Ett7cSveBznkg3OI4q/c/2+N+qC
NH+3RtxRm/Bh+7z4e6Swuab6mAmGWd6bTwJTeS1ne7fZMvYoloTcwh9kFNqasx2Qpq7GEjVIUV1f
11eBWZUdItiJprCMXT1+IbgfnVAkxqH1kU+qhr3qnoJcTWNb3K5bgbrbJZ48IRVi4Drl701ttAjQ
egs4/uDz/Q2mMFveYb2IVYMir/PFd/7UlB0JjE9cDzBP+3txULp9BXejUgkbPSloHFsITm/xPpjK
5jWsCQud3B+eDdmvGWGdY86Ume4gOiNk3y1ZUBOudwkpfCkL3mgBBSlHEQz6mUoa8ao4TDjq/xYO
vqSQo9cS7HiqvWV6wjsCn+zL6DwJvN7aEZoY2KEXIhQI5/Fp15pHE5ct0GCLdaQTh21RpkfwktVR
DEBhST7Fsi7WnE3A7To0ThX3wS+JuyYcPUzg/gC1nWFJbQaLKiEmr2XEwwMLMMldwJYSEvh1eDq8
FEVkUYJyJ4bABdd7gaKefUnF8OAsGN65cWVakj/vB9fNKQpsOMtE3RFMoQ7EhwRMdC6BHC55/RFK
yeq9sRXnv5HMLNOq8hyYJVdnGobEZ650fj0D4eIcJGezaBx405RN24UVH6TxzD9loNC0NzQV5UlC
bHnvTOb6bMu16w+nhApfYBYClvrfkOoX+XLhiWp0oSDHnTL1DbsPcepzIwRgUY8NZVcPYSl5aEBX
ycF2X1eZlMd7AAyWz+gm8UCydiimp3ZyO7GR1jnewoYdmotfu6oYzBHtOn9MsnvaAqMEZljiBsCu
CwKl7w/hGAYcH3TSYHv9QpyVSm90pVQHC9OfoYMOfoMyQnIj0mon3E4xILOjNHq/0jDtl+gJW4f3
0wmG1Eh+LjwYNa2DpRwUoWB2gmlouYJJLG9GJaXjerxhBnBBDSp3d87f1ozC5JoEsycn5dSE5B47
eKGwJt2nu8skJADSXp+h8xS5UW37XMVhuWruO2bCjttuhOlzmVQ3OuUZQq/o6J/X65DCTjN0b2ue
UpeeROn6PMb6hq7v9NR8SUu4AzlR7iNBzrqob+pzJn3BgSMjGA/ztlC6hewBJStt3gKHaow63SkL
yRxfuiLwEroVdKpWyxdfaPGEyL9p5VrjNEHtrMzbIiBKqC2h0o42EUH0lf5XgDjYw/61GQDAUzZE
LHasyNIj30gsnUxLgPS9nrlxi9i5jMyWNKNmIod8P3Nq1OPZQNAv4jqsQyKTfspGMC5h5sTJOVMO
GlWdmggFj6GUdBN8XNFTDM+3L2yhpfsbPY8KpfGI5ZdWudaDTfji7/rPXPo0nUbv8y3EK5+a/i+Z
UjRGP208cMENzaM7x+qaYqJC7uOAUyGcaMd9pcaWyPgbV+PBsinA9OeB2pNH78uA1qBzOL7FLKZh
EoQiSqdH7rbV9y32VNHdVqprwj5gouuIV+YHUzHitiS3CuJukapWjxaCUi/IR9sSmPR9kMnTmqAE
igJF0jrbZFsEN6fwQM38wuF16YksttIACaM0COJGCDzOVk/UO5duvPwSDCDdVAS98jFN9X/DXxbw
mmX0VgUAYuHGIiORQqiT32j6XuzFv9S12NprStTM4n80EW9c0MYyfirjILXBtJPqAzyxaShvtdeU
zP6HGedRGkdccAmn+Esoof/rrBqvenQ2MhI9lOMpQ5sv8QqnDaJSmG3nGmsVKi2XCwO98floCWy9
zgxiA5EjLYaYwHi2kW93qw9xPbc/iHFOgjxwuSFjHa6AycidvoDwLRiUum1Z3sTZ9G46MpL9Pwhh
+EytL2nXvkEViVbOstGDfKUWpVMeNnOEd4IVUlgK1Tgcid3oKVh7u79BlVhWXBpmIqHD9MUAZJ1H
Cp0Q3WaZQNS2tPrtpMpm7fLtk/XTKsLlC7lEJ3rzA66MUK63cM2HxBB85cxzsgmgyHa9gk0jn+wF
/MFqPQmFVccmvaVsYmDpso7Ddr6WDKRh0vJaiSFFVsNKW8s9408LeacuuZsUcMEV0WxF+0xw00DL
5QXA6z1++LS0m8CEK3zO51yVE7AM0d3HdRCx71QoUfevxdGjjqUOBuMoGf/OxdBd1+uxr9PpzJOy
QgLStCD4vYzT4Dj5AGzcgFZnZiHleDS49xbSmkSmt4z6QSlxDE2db1C5MKmE0fepLT0ZtvaLs0gs
HbLD8dSmfc0C0e/sYwDKL1L61NWXLEIUqldieizbayUswnuNwQc7vs8YFBD66lhytKPTRvXEIwCW
bnD3xDlLBePpHlu9SAXvFAqhi9sTSkQRaF9BTtBdhMb2IetPmYPzk2ynVVgN0nq6BxlY1psJteJF
JLOSh3HFuWz9nO9C420xuC+vId76Yo/OVbr5kafbRuoQdTM6O4xTerSFDcwsx+pGTK0R3MhD2oqW
kFz8Z0QP3majXjcA2d6kQx9y63yeEblzpQBzFqH+N26crQ2pD3uDlbbcQzO18990CWTteKLaEM2j
lnUd/NZWDcUtp8WrWUSX1j01/Q9XrggAmt1jxmi3V/UNwArSWxvU53kPFsAgr/z7kpu0ghZ6DWFK
+DhOKn5bMUSXWcASqWhiLk793m1zJKLmiyOainOF87Ha78svoUo8ZH1EAgGheGaICWiUTuT6LPpc
dyNTeLF0ibGCLYv9IUK5tCGSORSGa5IOSu9lIAwJcGVArU8XiilLanF2dExxSB7V3KEoAR6iOZqj
GaFeJ5fAe46MogHiobEIh3X+B/VO1O94tQiNaH/dPZR1HLJJO5fjoK4Sfv0oERVsk/vHtvrrNcJB
744plWXAa/Bl5QcGSrrGcwE8wtf+AoI/ioEeLG1ywRqMfifWbqilsG/j76SzayVmepWqaunxN0e1
MG6zdOy4Y31MAvNyvWIY8fCJvZbLVi7wdY/eRc/c30ddzEVWuEzlDPR+DF8s0hkj9wQuv2koI6QW
jGlBIRh8M+Hy1O6S1AeJgTcFpG2Cl3K1BjXI5i/BUNB22BRVuvIFwxZMDMMRWAm2kHxCkMpoy8Rz
qlr1DLvZdhyisVaf/aGsVQyJ/+9thab/rO7S0db74FLSVoKm8OuKb6g15dmoWK8T5mileU9jaMyo
JOSeCC8m5xNd6Z910VPhN6xFDzWTRRRHGiqzAEThnChGrn/m17S7gFDTYlsVqFwFicfZ2yQE9H8l
nrZJSo7FXFdeh8DPivpTYRhJzqiWz9m7M/FBMlxl0aypdHhv9JBjDF/RD3oGRmYHFgucXGTjYXOz
IXcQVC5c3sTixQk2e+2a744ijxjcJTC7R4C7v/XvTIMXx+wUH+kPCL95A26u8MFjBpFIdVO8wsoW
H7vAFsHG3i3cq5qqGaPf117dIC620YbfB512mTRYR1QqR0aVPpZCTe39Y5zwy/zL2fCg+XXLAZ++
/s/xoCwfLZI5a668+zWqCUBG0PFpPrCVx2KnPRg7/iN6wHw7J2UTxreBTyyrcu4Uh7cNHnv5V+wZ
qLULrDNZEbNup0Z18qwcuCaTzuU+XbE7dxCyldmaHs2Pof1bIkGXahg9G3AqTHjlq0ka60nr1RlG
Mudd/cDO6owxjKxYGANhtE5oSig2/csfriTFVpyYbXR7PWk0qRAo2KPKuJjXWYMQcQzgYK75wSCv
8SUJitAfvX0dMTqaEr54xd1dCriN1H+pwK99n3Ee5AI+h5wO7CM13+RFiETH1av+FlEPHW/Aptur
6sejcpIY74PGBcyBwnePAeI67FWOp3u3VBojg8TU0NWOdB1KzMf+RHOSrd/KtqZyczNhJQiN9rEk
MDuK9nG79YQ/BG4HgiqT4N8wyqSJ5yXMBYf//EBLIyyFdFrTpHo0qdfX1AiQQyrcSwt7es8a2YBB
KzlLz/N7SdlGXKVLvzNZKZAECRWCHRbW+fcnkYlmS7HZfwj7YG8/AellsrS3aC/L+XEGaarRDJYz
1n+pJI/7PfhYeZQbYSmXyBnriCo0b+5G4giqgyNvfOsIFilDPowFGP59GhIPDunbbDkGYxxt/n72
V5DJbTBB+dc0i//w2IbBxm4GYFr5e/QDODdP085x2SZEqb73+sPqrgL2ut4BBs9yS+r3H8h7x/ES
k/49QKpB8aDNyOydN/HdSuy+kurOY/ki3eYJU2Fohwhfy9gw4R7opi2/S4jx7yJk6kNrvLaKfuLs
Tg/qaTUCohED/WeNtHZWgmfbGVL6EYF+oQ+xkq111S9KEBhXq0v25flKnCISpBBa29MQ0U7cNivC
gyPemh6BLzBEVsJ1FSpsR6KwCIpheefUV/HWYkUjR3lAAYvUdGAGRpQ/PUuoMXCVPS29CWlBRjXc
UCzc+RYskkHCpyOTBoseBrsDvI+QFvA+4NerrEmByscv9pxzs+QI5ReWqYZUKz++JQGWux7DecOD
BCEUiB+FhmDcOm4wU79qlHhkkKxH6n9D6p/UdCxJULick3FDZtwQ5Zw8bmxw4xNJA9vrYluUfLGF
FDcIob6XUEjjXgKGpzoVCt8D3cgF8HPfiAxWRW7IHFdYw8Dc70Rvc7dtugT0N5tD1xZVhWMmfGxv
96BMe7mpSc2YijUtAlsmdjnA2NbmWQ3EfylzSYcrLatqgRuaCXLCkqYN6pWOJXIgdBvgrUlJiksQ
dh2tTtjoHu6QIWUWPSxtCwdV4s6A7Kc1tmMgXB2gGxOiH4UOuoE/z4QUD01GPGePgw/uulj5ZiwN
x7xvXHeSg8kwAV4SSBU/bYUs6H5MWurSUxke5jb0CLGusYBTQ7lXBNCQ3blHrGh9PGVK2Lal6F7J
esBETt2xXtu9SjdGg6XTr/mftSU3fGUMQGJS5qzAFMWiVDh4yS0Ys01LsSrO46nFulH7EBKfI7cL
eBUgzpKUbCuXu/xfoVYjyPbO5RZXvWCREZ0Mwl0T+i2n6KYgXFkesqQdEMGaO9mY6NwdNmcoPNXh
K9w3NZfgy0nyt/EaRPPdKwJ2pzoASAo8iHoW/7OLl4NrAzGQONU4dFPUFxPEuTXW4gX+KxoOv4fy
3AucG0uCb66C9rFU2Iw6kZ3YWMUuOX8br2ksAI4vtrkl7+wwXX0Mx9gkrjKvnt9uS3oeGtv+8F5v
Niz3gIpZLZdHoJdObdVsgCZHHp5gzHwzZQ9nftYoV9FigC6mdLwWn+x1SgHwuwfCrTRAsLDTbegD
b7tosvYwd9TnMOqpfhTFqajg/4SJK5DiIgKy4xPiFd6PlcvibHkDPUMAIHnXychteNfcsw18wWqJ
McahPpZz2dRPlC2ADhhPS3bvCzbb+LgbZkWR+0dXdvaZGfQdwANWL0hbYLhjoeBFHvVn3OGhTQzo
P8uY/1otpfF0HMRahsxGhDKEM5fIdt8Bti1GWH/PXg8R1KZjNuv48n6W/NoXRUzmnsuzZ/krPmzp
H4csfBDn5CUrpEsUY0i8UJWprQiq+jAvdktVBKTY5riYEA46VYjMnGlNQBbjAJRUO4WS60yjfCX8
w5eTL/8TLnRAQY3R++e1kDKQaMx1i+1oN5P52QlB47jR4/PWEM2kck15gT5u1bk4NaFdM+5RGf8H
fwdYQf4F20bAin7O4oHiDOb4+90F57bCeYeY7/nJbbI/5Nis2uhVV/e36+zNEjP8ni5KlkbIVurJ
ssfa2wq0pLxuPn13UMpWXkKun1Qz9BUtjF9GfSzFWo3i1c9EKf2JcumW6+tzTHB4A4CvlE76CWde
V1qTiXU6+G7CaD9+tNtd2UKuAXi2Ek9UQX0Td6Wu6layHBw3cWRNnHpFOB0JKxJ53750eNrVDI4v
NWho3V8SvPf8TpgFb6caO9WZz9wDdiu1z3XSheodmBeYgoEOCi2FjgJDzZzuURKjRDOxO1UbP37+
B9aTlCTbnh55xb5bGi+wsgQcz2aLZCwduOQtRI1orkw8f5pUJSophTroiJd1/yuumGdf3WcX8rP1
59woXpBGE3W3U9ZnZ0QkEWXZiBwfHDW8hvoQZCyFkxv/GzIGvdo0UrAfHG5q/cd5GKH8evG4Yns9
DFwFhtSGB5qooSUA/8pOmN9vET0PdL7D7ByFxCnohzDa6UbCpr9EJnyFLvrKw4aol9oreGhuqNMo
bAWjfRLcnKNG43naO8NrN4q4Adq9DjZ/mJ17D7e46XMrMHEHenK4h4e85s3qwmjs7HGrK4wa/CyU
CO92p2zG9bCI2FhBXnoMfaT0Ysndb+9QKBeqm075yWVMP+V9GyRcn/CBY6kDCRvBBLS+Ekte/fOc
1OehfCzqPS5AJs/cAyDevnY3PdI21yU10NU/femredHbmg7uyTCE0zVAGu8Ja3xajSDlWRXmwTu4
Yh7Xtd7EfYtz0iVFpSdQk9WJ0fFPEQ3CMLHNN8L8js7JLy9ykJBIfiP9R3WZ//ferHCles384yVX
7yN537Yz9N10OryZiLKXyWDz7YaxNHQ2gWuTkm4V9joWY0GUL9hqs+DyFAfDWOSA9cZS/M3LE0++
+E5N5/z44DEZSbGPCEpRyjvNoLktvW0P2OEgA7/v08WRz6PgweuU59C6IRPuMODqQh/ZrZPl+uLh
K51bfhSQL5cHO5QXvNx3bR7xv0PVBqjsT4KMGVNJqc1WyER4ASfdCNzVHCtbVKjSUGP/1no7ogNx
XLwR8qrXrEEqxmU0mCk7YXH+FrrB0Ti94BMmfqLAWr4zMMBjHPX5JLocUpHLXA7WQAjBNLT8vIys
lpRcgRUksenweaajy3qExayU0wyhDb9VULIQ6KLoGK4w2qX2qTXDap2os7Ddpz7zMOq25tKHfkCI
U2GYfselfOyZ86CKEy3wbw0ztBC/vDkXgyMKJt7YROusDEb39xyJjHPXfMQDh+Hx+qc+B8C+G5Up
dUAEaVSO+iL5KXpIy0m32f6nAB8xRLYUagmTFR8kvSLfvq7g3S6aK2Byv6lRYt6SBmglEfMrjG2c
Wu89YXwPXFQotuIcghSKe+e/0Eq0RBkzHQWDczzTXCJo/kYYWfLc21JDSRqGaVIU4A50GObPi3xa
PVUYk6d/ypjXUt3z4LErDzmLLem+eJsvjaYrjFeFtOD2NG5ghyPzj4tzhFXxlTEzLoFWroRxE+aX
fMrTZ82QWrGqLjhVQSzDhmTo3v4XTp6HZelSMGujglc29UGfmFnl4XHykk8xhKz+jsD9HcMd6NEh
rm6wxXjySXeIgvcDAPhmKeUEgUAeq6VCyWo3w8Pz3I2BArzL3v5NUuIEvpjYWYdlo187G3NFwTNa
vN3vTQfwFM0glGnD/zkl1y+vlcgm8H6TcrU6/h5oCKb6KXYhymFDh/SVcD5UbENrQFeDOPEgjTL6
pBmrv/Q48Xp4QkL24QFPwGDUqrs3AAs8r7yyPhchKfNe4skc++MpEcrnFq+e7k6/8qpy2iw1skUe
U0U3MxOZ2zXSkpFsevxMVTicIukw7R4Rb71zyRqYim/ZIJnkrEwFayCgsq38EIuPpdwH1KPlZMbx
Kc0UeZoX86SIEZ+fGN1jRzbhVDff4LFaE8qgHL7QU51GHYbyR2s/JY8UHDvIwe0CAdQXlmi7OD0R
3PRMcYi4VS9EZJGontL7+3H7Hf1UVLKdQDVXvUCXOitu7Uky8KtqEdky0vjnpdnDN58LJOC6550x
v+IfNBf58cflpP35pa4jlU6FXlnNlQCbchE1m+a8c5wG5q00GlLtPtZGHvkxa2s0+cg+Pucfs9SI
T3O/QVrrL2icsQh9r8HaLGmmZuwEgbqTfnou/cyZX5wtxdqcYR1QpGZW4SVAWjjEqvqH7+8lMXVj
yi/K3vtHv+SuBLIqE77YhkMqogUZCDCP5+s5/luHK3URNkBW24fOgJJVzs6siGkXMMAz+Se1m07N
GpU8vLsfEL/QiMh3+xsVs2sUOb35f4PCIGlVNy/DWDlcrvgoMtdpx3hk1yss6FTzFI+FLdldcwDQ
QMigZ6Ux1IaNWP+K0w85+Yp3KIoxMXCJkYLydDxv0xZUD3fp7L+/R4weY7k9j39ZDwFO7mlboabs
oAVzUXiyZe/lKATzEdCov0cly4+m8PTzC2iCZAjrDQ/7iAQQlsQWCy4tqIUPgUftPF4BXfCqIoxd
6Hzgpuogn3fWFdhJ4njSQ3pw44VYS+6evpgDSEqLIHY0iJpkrVK2RAQIqjZIgEPx8M/m8lZ0yuoT
uqHR9+3qfZdLtxMHVWxoR3yyT0C0BgERXX5xzoR/+Bk/w32ePBDxusKXez7ogpicb/R+Cj6XGJ3T
L6K/pII4Ur1zYN/TU6EZPOSChvfGCVOnLZ08oZg5ubQYTO9gYz4CJS2PJYgFTpCQ4YYtO07zAvX2
/nR5C06Rx05aYdVc72zTROJboiWBQmEOLvHckJXKDzvY5e/Cy07pVuMvuCBKUm5AJv7Fr3ptNbOi
R3I7lfRXfv8U8DYavTTWyhGlXHqYS01iYb9Zhj4/kHBVf7ATZFZjjyo67Q6GI2g2FxtbddiJuRF5
TFcaI6UG3sM5sz2H9g/EdIVhIGQ7924YQC3900pGWigzZUP3GWJ27K8bRw+DkhnDZpr5p0gwDpqj
Pv6TZed0J4THBXCC91q0cuJWyBr5GLJlKiibrM7zqJhMIhHjJyGv5m10V4727SVkgJa5GnVoI9cO
MjrUlN1H1h5h7bExgPZ8pJaR0JE4sugEo+3nCEHfVnf/un5NheDqr3y8VIFlR3nC4MV80YP6wkXP
T+BRoHKXuS6m/84P6v+DaV69ITfqbVSwtn+ETndEjeGFxfuylhTWNQRwUZ2Cdj/1qUhYGOLW3uZo
x64GrJ051/UzhUiB70sovsQfy5KAOe8rVWkME8FU/JJZpHpxetsbv1874asw0FUjPyi3GbN7cVqT
0U1eW4Hc7mQZXB93/+aifny1pisrCy1cjLLM62cHXVydNS/qBmrZ3ma/3EVXgQGkFsOdlhyFjaWt
U0Ac1lfZDucfID9X/kgzS4w0jXQaBb1LI1SMfx2y64ciedpYuWx2UekQDLiH4wbQXFMQb3q+VCeT
giRGtzzMbYA4ALO6SIn9e/940jjv+1qJ+GnwHsdoYn5lgQYGDpqrr+bGz2tc8QmaDXze63hy5aX9
FxSVKnfQpZrKDb9Ly1xY9hUp09j3CRfEoExPr4KmZWoQ3E1whHwBDjxD0j7X+BFJWbIDW3ZY3Bj6
XQivL5Wx7XT1MvSSTOQIT3Cni5MXFsCr3qnMaUaPE6/atvrYEvK1n2UGroKYmFmyiYumuzhCNaCH
uk3sf0Hr3RLCcoxhbS7VzH9PomV7E5h6gGDy5nyxgZOKrEhWqDMyn/hBUfywcWC9uzo5A5T1EYsa
opPrveonH2JZtJf0KxsFSC+oHP7vY2zDk0G9rK2DoFqbWzucgAIRaUddCmtSTquX2x0OKjEuVeT+
DIU6ix1ZYZS1KjAwjb/LYQeSMA/RvllmxfABuXAZlSngOuWHvpSu629o/EtHw1E/6T5v/SCHTKcv
3Wy5+jMxUZZW1RTHLoev4eAckPZtNeESwA5qlIJfQPK2+mkz65CycfyDYbZohQo8lgbULnhGCzN6
CeRc+sjlr6Z251Z3Cv48TAWLgGHYcid9HXPlkikKQezhn/ma0FPAO/VkdLbxPIrnNuBAdMS4wHUg
KEPQ+P65jvb3x+5gY7rR/w7JL24Aqr20fnDEcJs4m2Is0dkYQB3AOvPtr9h+dQWgFEBKQJv9984q
CLqAbif03p4NKOhBZIqgnBbGXjFD4ygqEkWkGE9A1fjuI12dlqXxpecsBukbJOfnowJieQMelIp7
CuwUYpE3RruYZByYKKIIenjuEPbLqguiKzSlJFoIbCQKXTr9fQueLcyd53hUkGyGQeNuwEn+ETqd
BG+dGeAzW7bdKYkDcov8eyccPkCfy1ms2z+V0jk6jch4P5Xp8RXNSBsHlP4z6RtxYh2pJnIXaIQ8
5HwsJiEbH5Q55kWayPzjr6yFKGHl63BIYzX8lzD1nkZ93TNRGdQC8XCIxTScZgNNqvRMwpA4rGVn
wpZ0pt3n85oodTFmC9fDV4kYepTRvYzMN2cDi7apjYkj9lKFsP8o9ef8S3Pt76PTdpXtZQZqyISh
9D973GDEMHXF/BkbCIwJ4bGUxX82g79Iw2Ck9yJ1UkTm904SDe6yVStGABtMb+Dm7t3aXIX/GLcq
jL8RaeKB6PooRXcVIjA/TUHfk1lQLpsGxyDP03wZmQLjEQX8QkHvQMQaTulBQXRBuQsj39CZlibm
WPPEaha0pF9ENVQrmCtyVKxoU6WSufR4ifuDpadf7zI/kWM3YzC+GW7yvuin0PIPDbkJLDz+ywKD
aDZLGt/gB0NG+aC9ldFyV7eOH3E73+Ay0cDb+S/7fBb4jOWFn9PUA9GEE0QmwvRA7tNHOl7l45+9
YMzeeVOMywt7PQrGGKvy77yPYhK5uuaCF7OSPNHo3tubegc0bS+P711Gh/z6tsanmY5CNDSG1DOw
m26JvOLTrjCbrIokYqXblyvQ2GQnSHeHtq2F5EaOMd/awW3hluS0VdHwMAJvcCrRkK+DJEbob5QJ
+SGwrc97QBs28iJVsGsYmasTKWV2A8033qaSpxmWmq8ywFwyhAhbFT/+DMsbM+6yho7zq9/jYNOG
VDXF2DCjIjlfU58inWEM50ewmDgljoO/2mZGxfgANZU8afynrGwcJZKC64nPGQ+gBJ/S2boaqkZ6
oz/nT8OcTfgTo7zLzD9LRtpNmJYtAENbcDA/G1ZPapXNA00UQT2knCjo+C3BpjCpGugDnaJlZtgj
eFJKpel3A/ckbHIInfoIvoNCAjT+TRbByLbOy7+slHAV0K3/vQb0Ruh4FKcBkZXG2FTgrAebfGi3
W+v0lk+6YwKA9icOXk7g28BroyGFlsPlyYT+wiaqwb7ovul3Uhps+jGB4H+thfCHpU/nHdTO4npC
ePRRPrH9+d2Hjwx9IuRHINLyjdXuWO8gNIVjPdvLpYu2OwbKSeuuHVefyte1IIfMdbmP0qM4BGTr
wJRJ3jAHE/mtfBk9+tXzT+uP2hiSc+jMJSR/8dO8zAIzeygJ9xQq0Zbv49s5eJ33hYH4dzcZG6d2
lb/un4yjIYXVAkoAafG4N1jsls7N5KyBDu1KfTg7t13dfmN95OAm3XUNqBeMWElJ16aNuUApd6pu
pEhy3EFRzNH/rE+5/+6sjcBiAuHGYYp6A9SFq99Lz3wh4fOjfA7cwI/7+PRt5mKGzsZy3t/xEyMU
qbhgU+BO5WzEMG0vyBmo7aYCBXzuAvzsnrFo37H63hqrJtAEpo60rfKPmTEhKuZuPUHaxRsdkq+T
afpy7fUrd0WDB5wpD3qRLOCVKE/JfrsSmuL0m6EGKAZiSHNFxkQLgClOXodwaJpnzUAFt0ww63t5
3rwcVaWPBfAg+jTJmhTdhLorD+pAzyCSw0UOGaZJO48UMcMhjB+s8qT2qofWloz96eD08UELyK1+
hYUJ4BqSNvBvpqwX75pEDg8Y+20vYkGTYrnwJQDhshmGA+mn2d3I3mzHfA/DORqBiJ2VDbVHLoBr
6tVqtlQvan9Xf9yEnlwZ19xSOpEF3TlmAAsVBtapyZgAlwMEgVDqtIN11KGIMA7mHY577Wps58HX
08SJul9LghGZYfdpoSsQCSAjm3AKI7cwrN0pQTGY2EKnmYoD0okgiBK6dFDy+qPiDUp52kaemV/g
ZWS8a54w2wkdUI8xt18m51KKRrdirMDTB8mGiPIhD/Jdo8BXsVB15Da+RnBxOzdShTpn77Gp/ehz
CcIlSQB6q3FychSRCLXyQ1NIjMs3TjsuEQp+rreQzhYEXhRvwmi++L3wNw9dVOPvirDzgskvOrx2
qwah/aQiKLpOX69VahiQjk/XxLm6wN7H2OXN1r6UbRylx8yqGXo26EbeCatUJcHvHB5FppdJ7nZT
Z1qbmcBn26OXhgcEDW8bRkicUrUay2R9kTow6GgcN/HRE9/6hdFbWk0KpUp2wnfdux4HnHJ+XIVh
hATS337ps1+4vt65V5t6ef9BtwQ3nTKgk1SvgymPC40rACzXgpgP5M2RfKjylZZIGQp7+yl+QSGT
zQDajC6XbmTe8hcwlxsL55nRvEiDTMXktEOOg9qx0w/OY+eVYDpAsJP1gc/dI0CbNgMz9MM5yY90
VTn7EwxDmD5l9EgkFDa8pjvDiKQA7x9wFisqPUGt26kU3Qt6s4IxNgyYrcIHoyO9g20nuRt5s1wS
Fgnb1BXg00JBcs+hbA1fVNq1X8EYTjlmzaI20b+EckcoJI4IHJEZIerIvtMUwysGlywrnyzQDbRO
hK7WpsvDAwa6gS+3UOt57w/jV+LR3ys45iYlZlGKpXDexr9xgVsPPmhRgHjh1FWJgiocVy8KECA8
7GdEF0BNGGmwNXfer+3c5mZvZWxgf1049D/oUAxZuJaxzXcMNVqzV/KkWFUP76D0jg3SCbn2jbOH
22C+1LV2PSia9YKlKMpIo3OAYxGfs9OrMRifIoZ1+PpLSTrSWiLPYelhAOgxx0am5RRKvTtvGGT1
eSSAVS8UxHX1sT+aYUZtqwvFBZfQgeQTbKHSC20nEhTCejzKHn3iUmM0r+BMc6IEQWou3t447wkK
dIuddv1EXOTFlVwooi+qR2NV9z+MLTgfgPEpkimy/q4+YfKnIt/1IbI0atOyQoDEI8tgS+CdqKh6
WR+n2ufkhsLsVQ/ZV0RPLox8wYMonDKPF4HIhU4kkB57vKg8j3OEtq7XXIH7eFY6DCPwB5HVHgKE
vS4t5MokUIaSIfC9y+ECW+u5LzVt+PQMDNlc1vRafeXPz5Bu3X/emu3mxEuJL5z2Z7qJT79kyWLa
MQSFtShhum3VDrjHUdhFNdK7a9jThRkIP6Unm+6VRf8oVoROzkl/5qzylkT6N1/nHQsIsDzJTV+W
R4jDxz9oCSr2NtvL44TDmoDKUCgBjLMwFCCMXIhYTE7oouUDX45+XnnzLlVep37+zPYS9fP+cdKP
3dZW25GrHWBQaZeyQHU/i0mm7cjYZO+qVBocNLSAqjf9WRvyWKRfifrSsi/tvCI3f6Sof+e9k56U
OoSt+fJP/hZzYCLBrTrECKcwTcpMrZcN9Nuv3x4S55BNDXfd8H/Q3gXDX1HgndIYoeOQ5ZB9dfGJ
aZEdKx2pjLE2/TU8kBsa/O7f/QxRP9W17rrYkpYG/oEz1rd/o83HVy2HSE745sTiLZnqcEC3kFzX
vkJT69pXxcbAdPZkqv/Cynr+LB1pjXU8ufySPxkpzZJTXzBYjrzbOmtsPck0YNenq2FWwcXvwzZ0
l1ZGSuHMJXxCi4YCqLgxAizhGbaDhV+VE3WI1tUeG+EybKSPumaAibwIzsieszrYcDzwC7Ack1zZ
62/i8J6KvUgcFNHp4eKddtfnTLSjeqb6gLP5Z+jmfyuI3lkwAgRZJMwTMXtvufPanWG4BHwBUF8+
4Q/F1nETMIEK1SU3MbyM3ZH0mhXOel/DnHOOhRoYKcG0Vb/ANcpFhQ4JZzLmu50cAgzUZv/Ha2W6
pnOc76GZ0Sq+wbkah/uO65PIXFhQrqZfEUsPr3Nd4M+5OFX2Ho0+7KVzTHiLAqb7/ui6pmsl/peh
26CGIwmU3wweXrLG7NHgsMrVMfBadrpTIXZedtdspJru4symsQ2H7i3+LGVX5yeK7vKQEHBo92Jg
h3KXz9bgCtSAGJ9m9Vk5E133GBTwnAy4vcMdNFDfGxfCrbjR+q3OfEuKWAMl8BUAPXqw924Wm/X+
v+9JAAYFqVelxNoCMB1LN8hmnwKBVQyDdBlFksQNSQpCPy0H3Qr6lQN5Fw0tv+8WPKM4MR1B0lgC
8jOuj+pqywj+nJ0OdkEo+0QKP5Pb6kHR8wjGenRMBKmbt2E0RcYExY2zLjcSCMFvR3JmNPobl2ST
8rcnKNhOVlabKrDIB1bgcBitZCRSWsrhoZZxnNOEYFllK6JQcw5OrWzcsZgwnOdq9uNuoxj4x9CT
HqzAgSJDOyFputwR83BLH9ea6cg6mNHNL3aKCU737tl+foQaUf9Xmcc7o0HplS1DYfbxgHy4Ybl3
j5hVQ8fABl9LQYOmY/XKFoldKvuF8m4yMuy0pnLFSJ4Qxc3L4L8mfE6ukExCbaoUT3kVdDpeczQN
uI71y4a+trUyxk7bHvq6t0LZGhGwhNYHQUAUK2W2FezZ1Edx1bcmVI4Dni07DZ0c1LR0oZKaeZrh
lrsJFULnDjEqXy+8Kpsorw3skfe+YknotWFat4ILUfjnwJEYxxqKrfHXAtVXd/vKTvDcWFzsCbMu
s9oWdr6ZyHNUlxeu6tq2kRF/M1Trzp3b9YRhXCCCWwtS/I7smb17c/AQ9rWWShDTHA8Aor7aXDcP
tKeIYEyYFXLUBKiLclLbqjrZIekTrv7anOURcEqLQtz+8E1Uw9u8L09YlY2TT56QrzWuYK9vNXZG
bWcl/40OQOLw6XkcVSCWRRfPraFUWnmFHNDZKZETjxY/fTcvxRIE/Kmezot5eDxtXFu9wAoB7RKw
X5rolZeSBMeAZjv3eYYj6xKaAUqa4n0l267iFEQDz8M3c9rMOIWQho3BmUgC0/sp3cfViadyLnMr
q2YUNCKOnggcwBgVnTMSMAnpPqUSHQvNqI5lLXqoUKoMgyYChXrfxL+gTSScy8X+ILJwcuMHVkn5
T9RJMNqsmG98unvnCcArvCkvYWs8O/9kTPpzxVHpcG+MTNwEAjwgfyXlViql+dlhPoouvPXSNw1W
yKJchZTPIwQusyTpfDGNT+F1i/txakTpFcMmPBWJkmShMUFRZ0oTq6Q6R+yc2pKshxe8t8nZshXD
aQW+Nvw3UyuCn5CxUSLuZgfsFMOTHQEVJG8tKbTO4IvmAhkhOYTJmgIiDCE7hnsUrcnGW5vGMz/9
/QxQJxKWNTJWr+j6aRw95jPMAA+WSVH1uxOwemji5PMA8L+Rpx02aIc06Ag8dRMXXo1wk0AFl7EW
zrkzqv+0QOOBz0hUMzZNUbBbVy6ZGYCMnv0fm1rBW9l/h7SSsaC1Hf6oeSva9MNOU6msQBaKfUh1
P5iweufJqsTVipiC1BYWQHquD0q4tmoMX2wHmNts7lthX0JOmZNlxHsY/CF5qwBv1vfqsO8xHmCk
hwNvp+NWVFl/h2pk/LdNkfWZB9dXMRyeIOSA5qMnnx419VIAnyF6M/irt12jnSTNFQU4oc6uEROe
RRYNlPz40VFwR8Ds4cMNfSBmfHIOOhzKyRSwiKtmMEHMX6C2/JRg53f9514woM3MJWxaNd+CJKAY
AdNL16+aoX4rzkTQ3vGUEwi4mMId1F7NkI9MNEOyKfpPT9YhUnh6cq8swbQ1DM6QVjTw2cKY8VYf
zFHiTknEMT1GB9xRURw0ZVYJVNvjslU5cbfia33WDppv3R1b+L8nIPXmomI5eEvVzqjfgI8Wkz6E
uki8d0u26rF3rvT7MGq6AtcUAEsvIbNFvoxNEM8kBGR5Pstgf8WJ3Fkvf71zQMCWyI/K/pULIIzN
rm8UVGOhO2okZ+krWafOfG1qkVN7n4Ra5AvnoSVwaVCdbwcMRk1PLOzYFTq2G40Ypk0WulDKRdt0
N+tQL7YzrMQBMRpaXEa56zH3fDy3LuA6aPGp50OmNxCtXujFbNC/oQqvIZ3cxIySDggk5NFRK5k3
jqKiITSDhHQu+zOIh2oUaSo4rzLVEQ77kLGkZcambkJX95kMQx/r0chceiPKFmwmnaXcDuLV/M22
x2IHx35T0GqW3Sa40hUdNpFyY3ftskOIewLcfi4HAOK9wOB61PqI45iltPUwvpVY7fxo4cnA+iih
s3JU/Ie0JK1XAAmsI3D+11LFI8H/0hULAMPsbOzcHb/cyLT5Y8EfaWU3T87KjwdwtyVcqMRArFas
Nv2DMEah1sSKqHOaRNmvpBjcJe0mD1UwxQ+KCrI3d5tIuVAx87fCR6cxMeBfhP+XcsqT6GQ+2bC3
f/z04lG6FWEHIaUNxKPbUUQdY8SUIZS/E70I903FKNVOrNOlkkeaqKEaUWGWJf56k3E3mrloc5gJ
KgcEG23pt5fb2U/mnuTrjmO2i0zsysh4lovPA5aEzr6uyZWVx2DAkQM2ROKurWQbC0tvpLXHlgtJ
z4oHmsB2LgpXls0dK/UrCkPBd5/uG61Wk8Yo1JUw7Djp/V5JyhZXPWiKqkedw1mXD+MjttYnt8TH
iTYvzj6qqj9/pfXg4hzyLe43nC1oVOcP8DpZd5qgR1mSbyrr1jh3GFKvLpk1/uQ5N7HsApvoBjiq
o/3qeCpTJ89fWBMlYx+2bti22Emso8EebID/vD41L9qqg4Ivq0g4AhXBmERtD0Tlzzix3DHcel36
TyV2ruki1KRvpUBxMadVArZpNwxwZD7fDApglAnqP/SVNn2SJMMBoL+tV5KqpjTFM1b2D+r7EgyO
EKTxORDWZry1S9IsKUqQ3zy48T/iBbHDw9mfEPJi6OTQzUmISgEafqI4y/lbMXcYo8WFaVJCjA9N
6/XG/LJ9y6WuffejQFzPZGA5mOT8UA4WeN/T6ZJ/ShBcpui84Rirp8E5gIoQPnjv3u6Y2++2+rof
ihnawSJhbqI7DeWnrBH7tRvZup11MBn1OtS663pY7vqMpii83TQwa7OSbczFMfn0vJTtr2hA4NQx
5slbUaSjRtA8Rm2E+b18y3KL+xlwIaIl05ft+J2E3uB2uyGQHQGzAZJOWYipujTUjliJ7yvKpMo1
IKM+jyCr/hGhwpuF0xxOFuuPeE7JnLN6YgtFHJRLp/FR58IkRxYAWEI5pQ4SgyEVToX9Km7iDqY6
AKGc2Vw5xNxcVy7HYKL8C2DnkNV8Vw0ODCRgr4hbmz1CqM59hTwQMLjAAum7U/7cPMrAaCh8q2rW
0zjHTKklStAu59PApUTmSm3+se096swNPAK3s90R0nJaxsLUbr7u/BU7PnKA63qOpHsuX1eSB8kE
fEcW0WRkwj8R64jtywagBd0UDr0zihupCaC9gZS7ZW3nz9sQ4DFcdkFJWbRPf7HsAsLZSVcWKp8a
SFvwWZuZrxu6UMp770p0P96WlWtMjXoBWA0DgZ+k5Zopkfy+2bAB6UNoOgkKSK1AV+S7+F1nJgTy
mpxA7Wvs5ekOBB4Qn3mImy51JlCBvnMMeLHnZcptuhhGeovJ1G6zBwnRuEtybHiG1AKVgi9eZkkr
PR1txurhVuOdEtkiyDzqOEIo/XpgdPAj5VteRyJTK2XXDJFw8rLaDdkQyBXxPaPObaLJfHA+z6c+
iR5ymkIbrlXFX9uu/E3Z21ouQQLPGn4+Wsd0MZ2DgJVxB0h2u3moC8dx0ZF2u1m748cqImlPUvFn
pZoLNKL18Ilx7noBDGtuNhGGQP7OAfF9vpo6H8dVJvSH3bPJDI8+Si4Tel7CzwBr02RhqiBXGvSE
8iLv1vHo+NPGTsiusJ1Xz6kLamIWHFfjUZeDjHMLw3bTs4CHacB3F6h49lJ+fiuCeQcOnblqiF6I
Fr5YvSkpkYLWbITfTjPO3SGC/YmP5IPQ/+cdhI52vUd7XtkGl4/BDejMoHgTcjP2cZsbICEoc2hj
9l1iKqMInCRMr9EBIZ5iAUvT0Hspg2om+ItcyQh91qdzTLltjhpWEU57fnOawRJpI8ylocZe2E6t
lWFNuvd+5TUoH8cLKV2z9J527K5oFbv8jPvnWFw/b3MxevwVvvALPiahNmdTA2gjE2e+gLVPnYQz
eH07wZI7+M08lk/GMoovS6d+8Y9n+AH2rrIJrG+qBzbAIUqVOG5S4nBRWQbCsqJXJHEt+hF+etMj
SKaHgS0yD2HhS/drpbkT2iX2vEFmcJSXwPXOdpwUka258QE9YSkLU//wWKXoTGeajiMyNDAotSxB
XDMVb4gddtMg7H6OpWQF+ZDBysNIsN1avSuFrm+RvFM5aMESvcQnEJBPVoxRgP/m3unTdlMLSBWO
ahmbZ8tGIjCh/YXkOa4Y6COqt6abQ4+hzCzdgcvYl3fUNgQtaZ0H/bcZrihmkVlpj+Nw5D7hfXBZ
1xrTwawvbdM6EGP8HuZTN/qDi9VFxG512s6J82A8mhgQR6hQ31R51GvJapkRaGp0tcoSZjpyV0z1
kLtCBaC1hSvj+87TbJ2slfIBqNUHi+pv72tf7KVkat1vEUarzHD3Pb064tKYLHYetKEelwD+ceDm
uJlLOw48JCNy62mI0e3onPLdNepeQI73sHP2gANxn7fZ7sVcNEHDr+irt6WAys/iIlZBhiMtTeKf
qFbxg7blk07nJeblOL65NHJsqjosvMWo9oHegTp8+CrJDYZD148n+cqOB3zJgf7CgJY1pjJJJ0+L
TXIZEzbfNEib/Pbiw2/75lwi6zLxoP7pcHIBoJycfc99PAKk2kdiEpDl0Fyrg3uVU3bY3oTrI1hw
4ycJ+PFdyp3r3lGqNUKvKGq50NTrrLEq0LLUKQDszmb4F7JHw11lAygkL6I1Ys/WNEnlUHE1c1kK
/FNYJcWcUxxhRsi7XscbufPkkJ80GhtiGGAhsnlsU6UYvjiHY3Hn1fynd8OoqC/67r9SsfvsJzrk
mxYmiKOLF11sUrr6/bW5lAof86YYNquGx5TlLKCqEe4wRkDZccuGQBYSpGytw4N4EUfSVaER6W6B
/WinFPkDrHqRgoQ30LlVXhLA9s3MHnzxZ2MY8ytzdbr59GJx1pyoTUlZxE1IYPIjFpdY4d86DHao
jsdSJ2K3+VMdLpojVAafOvQVlo2npocmOom9Ee7s+41MrBZyEWM7leHfV6JzmSQL+QfXbIi1kJQW
otYT+icP0ZABUDUMN2nS6QPHv1GB1gP9iUGlTB3r77tIcWmuZD4XFE0FbO+5teP/eU1bO9tueDWq
5afh679zXQKxYVLSm5BYkwdE2vNcuX+HkrB3ha4m3qU3yXwIEPb3aGJoOhk8bCWIptypGv+6suMl
WjvFi5PcCZBIIvxU1f/e4vXVbRIfNk+twGr9iOY0t/RXBV6wD7VWdTz68j3Kp7/NYQUekKeEJ1NK
bDMPlrPhuleWvYzUe30bPiM8CpjkM1PZUxW8Q7A6VpBrf4zaEREULaV6o8MqoMNwC6VvWgVBTNFT
816Wt1glzAQJyY836OOESgaIOI5bNtEQciG5agMA96COCtswZb3HbvhZ1r79v7NIePYUDNYdUBgy
xtEJvZqz8lapQPbhJcAjNxvrvYX5Q8mOMy3YqpqiTNb+Qtyj1MP3LaW3ZkT3jwwpjvl60V4bDsZ7
UXSoSCJbuxhL3O2+wygTfqN4GMnCmdl0by6Je4E3fw9NnHlMQe0iv/kcwA/84nGaR28c4LJnFjTr
3pI5HopOc+iXEfM2ELrawl0F1+FpUjePZD5ZYDjOsE5Bm7PdQOYE9DQtfE88YAoDYMiAdoTlI+rD
RPEYeyVJm02zBJNKmYss0S0KZ70gd4si5kM3jlLKU0QkdMtjeQPhDuEvMuxiPy+yKFj9a0bZOwDO
gxTgVdXmVOK64aktPuacOZkOUAO6HPzH5+pZcP5yuenCamYcdY8gxoatj1et3MJTeBQpEhy2bXkC
bx6jTAwC3BNcv8CRHV8FIl1v/amdswi31rZPaFFiFHIKvo+SO6MA7nxw5mNP0s0O7fE6cjM61/+2
DPc/5hCe6K5xljXtGe+4jL+OyU8PuZLGPrK5rPZqcBDSHup0iydKWOCnJ2tdDmsyOqjJhEP3j+R0
GrkDCeTd5i47CDClho3J8e2Sy4OPewVqh8fB0Ua8cWQjA3UIW/LkIru/Y10F/b38aix9OVNBUAld
6DEoqE9koZz2qnT5GVCrwfX2Mx9soYSdwaO3rYt4LW6T6DHGClkBmRWKprieDYu72wVGsGWwgkCa
T1T/E78y6n+ENmJOZ7xSXJ7tSEl7naJuAc4dVb/Ai1HuaJpj3hzUkpHgTY38/F1CTR2GQfixt085
fhSAmd93s/Zw2rsJb9HFag==
`protect end_protected
