-- (C) 2001-2016 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
KIjsjm1OH1T8WPfd+J4p+WqNEzQZUsUPzGQbCfMKgzcKW9Or1Zn9tT6642IO9t2zZYn9rPcG0eZh
qqSeFZ7AqMPqH5LyQ+KnCveF0mQIClpwf46+EdlVSKVxgPysMbN8SWSh1DfGLFrdCNehGnkOC37W
8QUS34eL+rrku1LG7htm94OuHnPJLjEsucgTUCljB4Iy6g5QAoHlNmHAYaH0mVn1dFoQceFsNlQY
AbYZMsyV+eZzDlA/QFVMTrZMSwrZ2UE5zB9LF9EBYFMw22p+KrSQ7J4AYua2bVxGnK1U4i0050MD
TcfheOf9CXSatsAm5LiMv4oCsT0QD0H5r0JEOQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 3440)
`protect data_block
2R/i/PZ8Doqx+Qz8JtKNP4cLfEnmd+llBvcyxkzI2t9foP4uKTeeHWAG8AUmUG8WiF9GGgI75Mz2
Pn7yaYmH8Dp5HmtiLuJTpmukAEeoF4RoxIPpaTBTwzS528Wk2XBzAWCPI/dM0IIOj3k/XR7yArMA
GdFdyyvYZQ/uFOFIGuYgYkwBSHPDJ5lhRKotPdpLDYmtx+MI4YdkdxVexKMWZ9LcyftBwxXui0nH
WqplGQTTJksY4ZzwiMwZOuUu2Qme3jOBxSi+Hy0aV9pbVcRi8+8RZJ0ua5srNJsbvvoj7j8pWLCX
PdSs/Eu1j7Ko32S0x0o2wVDe88WdrHF3kqiIqjoUh/W+xCq9OX/xIuuLu4jiTw93YuR+HSF3YejP
yhMz1yAItS2mbwmQcb7EW0foYYBvKoiMcQbFtdrkbMbx7SBGb/88xhRt0mWvcC30s6DPy+oazpx7
VccjQE5jtbr3y+hDmu81ANxqzVOIb+uWq17B0yYGt8CZxFdsX3lrwYSU9KY7Wolv+xG2xb89vr+C
1/mfeSSWVyYZUZUf/Xj33bswqWJiB9rKFDL7yjoy6pfgrjNcldpm21f2662pckq7DaR3whAMU5LB
0DQjsQFKtplPRx2gPKVAmZZP9l+wPTqLeb1RJwJnBABc1KDwvUf8Wj9W/E0WxylEMcEI0cZZUnLP
B0L/yXQv36yWsUNbF51wVKjuKpxbrtNFlb8t4TxDcXJFIqX9Et91BM5S8iqN3wI1DK9tJFO36nNs
tyRXQnnNWzjW/4D4LKy421ueBTf667qmOXeJ42BzvX8lz3TE/XgpKZppl5maFL1P0FhDKb7jFfG7
25g47IKvNmajidxMt7KxaKRRkVBjdNM5113GXUlpghB91BDF0ewuV5gJiiRwy/oBq/rdmSAiTkwL
gGmIxlmtpPQsPTGCYGlwYW44agKexgz7BSoi7/7/NYO2kg0598uJuKRhzLcn6RTqrCzwH8u1ZGf+
ecJXJUM3oHluTVfKfH0UfuH9bKubh44lmKHr1Pk5rBrheyFrFYiE/Hg6O5vRDJcyUMBGcanBo2lj
8qowSbqBsij4Ac9Nw7Asr+OAHYVSiIh1MJc2IRaSR7RP74VFy//6QkcrXIK51cqw9Rh1C3kve32p
hTmT27FNXiYWurr8ap1yNc8/wS0ZXYvCnTB8Sx2nXZiKCToZA5t4rgbGS2fX9ebIurU9lovNOFTe
BMOAx2L/AZf+trDxSWO+YgirVWk5xJpeSe534xLpUWaRNadlER70idukIPNJ25OaXxGrXGxJsjbO
ReYJfQIvQ9sSrlWyAE7EhL21C25UHPEVpMAz3xcC7GRVHOc+qtj2enYL6dEzlAezaic8tnaUOnhq
7d47PUSuQ9k2o+W36VQUoLM2lL5iPYImh5LCJOAeMKATCzRoZW9OyJmH+OMIyI1UQFIvuKe7WQQ2
nlRNSLeyd7k+z+XIxjn4Ix3HLR6qWGm8/Bzq9ayV3X7XDqZZvsXNWsjPClboXqgGVXpMQLTSYFFh
4JUFSmWrnHOkDmU9IVOQNlFHG+wbXjkjNppJL5Llamvf5pfgkI3FLnpTXuvH9JQsTpZI5oRg8yzZ
n7LRkA/zSBNGHngL8/+2RF+l4e+vxzFPqUZ8h36vGhSjGvxJtfu63FJ5XYxIb0CgEjYJ5NHjdWvK
2vLFzJXffbusP9peFdfh60AeXzZ7ghrDyfCMgFyRFF+mg2iGLXyn8C8W4Dp2JFUDB1PrrlUQaxRh
KQsiyjTjMiQMn8VQbXSeC4sOWJ74jTBe6tDsOlv6B4OETAr+lS1QlOv0zENC9mKmPPweBNzGzDJR
uJDvbPLgr/LWuq8V4PaVeLV0FgBd2z+006Zh9BMFlOKXowN7w304i5tIg+mar+xLYNFYCizS2occ
h4IMLdqe7PCWbHlk8ODFL8Sp0yTYbR8XeaEzjBwqwsteeqZ4oS7TMLjayEstQhiI4XQAt6WnSmxQ
FeXfTf+JlEAaUtAbMRfRZpYKrHpaOhRO1VPAWoKp4fUCp4LGCobZav2EDrneo+IFUGR5a64jvOqd
PthaI2GLshkQMd+AM/aQvh0Z751aamlIXL2+YjwYhK2LPq9I4eQ/mHGiv5tZgK6MD/pYQ07qQbo3
HmJKrRpvtqWVIRwhGDfBsh2Ylww0kCseqy1K1ucCjwzVTIu5d1QABT3ruwDDd0ZuLwUOwrwplhuP
kVhE36hNUWibPR17jxk8gL4ZzM3hYBTufuQYIFyaINeVo6CPP6+7KLIMupXrfDriokWVDbZWu1Ha
jDZlB0mrFZr1igekx79X+qYRnRcZ6RbL3VTOPJBvthfzCbNE2g0SkzcTjzo5eZ1JG+2qBcUnMIPt
vGIWjDfwgW0otAWWgMTkB1UPn/M68ahKRkg442V0mJtnqFbF/tToj9lyFdiF5DTC+9u+Jmrohhsj
hAKtivPetyTzJFXoty2VyixnQ+qMLdhhJF1/UjnpHyPqqARgv74Uflt0TeCNooqC3uFX74gEEU05
Kkg5RiLczbMa9zc2NdffSFFc7XYN5r6JMmoC9LOwI6sqO9aVFARnIypIQN4iT/2UfKDqqZwz2CJF
+T1zPuWFTkty+RXvpxRB+rrvUfsB5ic1PWjFRE/JY49czphJhQECPiE44tb4EAs2TuGms8Gth3O7
wRf7kDD5t+E/lnOfqs9hkIxipEFFUFVro36akJviwSlsCcYS40a+uDyOPptTy77NpV4xq7jwFl85
DBJP0UjRzsJO1gHprey5K329cWtr+jWpo5suTitYHRfTouJImiQRc4zbfjDSrCjmc8F7bzkEbzCP
hxunJv8ad4uL4ZNqhs/PX46ECYPs+wgn21KZkQageyN0fxQfE8YlMLlHtyjrqzNz7JKK6nTPn7cL
L7CkTDBYu65dk+NrQuhEqAVLzCw+nQQ9o419WsqpKnnr7DB+q45l9ms1vND2N7V64Hio+Wuh3Iww
0NWzfqF0G/yzMhy1Kzaep5nk+ej70uHX/A6mdh6BPllamcA+FN+EVVcZv9fhfWNTKxee964h67tt
+zKMUWMOLW5zstw17tndyGFqXKYmU2a0I4VP5Lj797Jx83uWCeJBatsrjclJNlbFhrmsxDiufdr3
vc3CQX010+Qk4ebEmTI6m1j1Vr7Ox9xt/nyslvoOVIMimpw9a7yl7qU7zsdEXXGHxDy44iVMGyiz
2jEYIpK4KNNPQ8Ttv1XhHX/uNDCnEuzSDsATN3QvUQNJtTEVJAdJgIJO+i83NLYqBYU+FzOY/Nfo
1kiigpfZNB99T0H5PRPzwQrwF3rGVcgsDig9l3l+E9Bblpl5/Mi6hmZRnSQMhofzrN/jQxRtCe5J
5pOsPsKYFOn+5bm8qjHANPzJVIc+GZ1xJtKORWVRqURhqKBFksiSS0IidVgZx439SyD8EsEDXUD/
Mz9rntbe8aLZh/c0/K+ahi9Sk57cfEJLqfVbZuJEcn+uMqRx78d2iNLPqYbjTYU1Y4ivsdlFXt/J
WOzQhEvUG9OP2JgiQFx8XI6MFPsF+dJ6E3s0vGq9VX0mWpiGVTPi4QIHyoqAX+0yoWx2tuWF3SMU
o0OneBQxbHig5z3aEVFOoXkKWBRiYc8EzmngUh71O0GxSlg4QOVTraerhfTLOJVtgX/SYIlhrD/a
hv8WpQncCSFrpOAz8aeaKAXPGFeGRnZulyQRkNeKnHFLtXbihdXSMWan0t4b83zMz7kJ6hJk4pAo
VW+gxLqPnSC7zyHuXxadlt63CsmGkPPAvbOSmE1j+aNIMDP17z7mSJC2Do6gDsSYoazv0Jdo/OpE
LNfCF/0aZLdSsbH+F7FWfoB44FOIGW4A7lQItEOcZM1BUA0/btrcug2pzWjxs9fKXQw9n3eB713/
CvhbiAYt7AmtF9FFMhLLIYICop7xadc12ieQvyQvz+9avd2EAJWfV6DnT5eO2KoYJvJ8NMTGbXyF
s4A86gIc/bLjzB611WcUL7GHQx7xiwbCcW7ODVjF99pwVy3P0uaPL/q5GkTNZHucbirzwOaaQWKQ
8dOR2hISq5nkiR64qIb3RNeNrNyQklkJa4InxzUca4kpYs1gJEnWCGJtSmI5z/4KkeEe9TJDifNy
2VhPpQe+hE+HakQkoaH0EUbfn87b+lQnb8FuPYyLUolPr0OSgG5C4oNbEmgHF70ZlYJtweRIr9lt
9flMcBaC3fOdvjujPqH/WrTPMjfSYdN+ffkgvE1h6TAmvuiLBDGz/PHzoiPymvl1pt23ODjqTay1
/t0IPveLE3yag+DerzjryVNIt6qspf4t9Se2SxaCFESlxC30MFynieVI6Z2zVyMsMxCZyWt0Pcti
MHJlh3FY0ejSl9GZvZe0b6h3CxHxCgm517V/kokrCWkKVPfPQbiH+hBMq9GMRz6PSOAGYa/yMF5M
WfRBEvqow4iXAPS2RI1yeASdVDOgJJdldJzVFlFA6X9jBjelOlj93r0T8vk7J8UD20b6Em9VALbl
SMTdc1gx98jujuhkH5ZpldtVXl8nVujP4ml7lnWjg997Ig1tYhLk9w4q3q1IjEsMKBTP+jhHfZWN
2cTEHposHBTMmY7B+12Es/DPnbE=
`protect end_protected
