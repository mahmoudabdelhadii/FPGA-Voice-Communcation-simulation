��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���/�����Cc��<Nb��.�x{�>��0����=�����=8RLG�h+OLزV����ݗ�@��&�K��4cbXu�6@A��?��I�=��O�s=���
�S�i\��D���d3�q	��9/�I�w`W?ދ�S"K7��5�,l��C���
@E=D��!
����荾Z�V�h��c,Dt��&�����]4w9K_9O�=l�uE�w����[R�\�zÚ�-J�$����åCj�[�
����T=���K���h�����,������#�z~��?�G���B�~֨1)��k��yq�$/ju�YA9��SX�{@��mWt������w�F��r���������O)�mC�&�����$��^_��|�����=������A���_"�s���50��-�ݡ��kVE~�cu��'Ah%�����v2ݲK:|�g���7/��=Q�u�~��qC���
qSa�a�n�m(�]�h-�FK�]�Z<��K�b�s��'�����C$Yכֿ��h|�[@lXJ�*Qm?�аR��(�v�vlr�j)ڦ��0p�s�bv��jy�-����(��N�vהS��Y�n)!��\|9��;#�o:�#��9|TWL��L2=�'���$ƫ���19�?�:H�A���T秧���,rJ$�p}�a�ڡ�rn#9���~�1e�[e���!������{�T�7���O�z�������쉎�<o�j��D�7��lS�ƃ���F�V�:¦?�,�:4I~P�o6����2
�ԫ�#��G롔�qH���'> x������>I�nN1.�yφ�V�ǹW�)��	�3���k��c�Rw�buRA�8����\��L+pȓ ť�;h�%�bT��к�c&�k��+�����G�#l#̷ʥ��ڄ��ѷ�T�b�4��׭2���@�"RV~���k'���	��v�.���3��i�'B��3�;�{>�'��O�,ꈕu��醁�7�G��6�%���Ķ���r���
�0';��J�.Cд�Cz��M�'��«o&���sλ��˩�8t���CF
|�x�@⨂�PE��8M�0��x�r�=,�l���$=�֟J����ē�/ +�>Q/u.����J�o���i����9-̄�m�fEm��K�ʒش\��+S�<c)R$���Z� %ښ>��I/j�5"u�W��*4���SA/�ֹu�=�J�{m��w�t�J���U2�������or(׃(`�M۟� �l���4{W{��SЙ.�|�*l���5�̹O5�736J����Â֋z�h+R��Y���/9*?�)��ڭ���ҕ��ڌ�n�3��U�~��o�ܘ7����� K�?t�2D}��s�E��R��g[��En���ػ ���h�a��h�!v�,F�+ ���^z<暥V��-
Ү�|�	i�����>�sZH+�6hkQn�Vϱ�?"��IsǓ�EB�{vm�3���N�/��X�k52����ۦj���)���bj��54��.'l�!�zd@}�����epo��Pt�HL���Á���%A���4m�H3%Tz��k��I	�WTx/�<o��|Z��W7K/�M=e�ʅ�X��\�6d���QEy��)�˿Zx��Nt*I��Ha�4��48� Ҧ����ҁ�\R�Z���8%��ׅ�~S�i����3�wr�~�e(��ÃpȚ4Nɼ�uڢK�8gKX��e�J1�2Xv|l�+�ƜWY(�~�<4D�-�aI�G�)�!]�K	y�!S�@j�}&����$2p��ԋ�{��3Q^H��a�S�(�T7䶡�͕����hIW����O��nWC��d�%z�R����Z|;,�����,o��')�/,n�+���]o#YZ�����c��am�	}�����2H��˂Zk�7p@uY��u�?f;/��z����4��xK�޷OԎ�	陪�CR?�	���i�\t ��y�:�h��.^u2��]���6��BV�N�E�G%C�yF�E5?�RW��FN���K/�\,N��5�S]3��f+� Q�ac�� H��%k�����}R'N6B�ᗐx9lG��ȭ�n�S��>�s\C���K��'X��Q��}�v��ZI42h�DЭ���M��	�����\t0XE�)r�7Ց�����H{Ҡ<:
��Rɚ("Ð�f���;�]�=#R���x#^
�ω��^�z����7���A������c��J��|@�;W�Y$]t��Z�JW}�A�v�%�/D4m�+*,yu=����^
���y�4m-Ǫ��Oi�=*�U��?�;��)�Q���89#�1�or4+�b���X� ���\Y����~@��@v�Qh�Ԃ��D$�Xk�0�F��5���2hǣ��C]���ס�`�H��ܜ��I^���\
S�M�G)R���'�2���L���*BռC�.��v��}�zR+�* �0~)���&=�~�������`�RTm�f�~���-n���)#�������)�a5KU��Z%�3�l���| h��}I%�	�J�'ŉH��Р��ϒc��(�^f^C\z�|T�"�l=�zIP�{slͦ����١ڲ��I'dI��>���x�TV%�>���p��)�FL��گ6Qo۶&�M�;�M����%:	��M���b�5������+��%�Ęl�i��f���/� y[ێh#T������Y��[���v�����Ny���!SO|;k�k���;�3������y�X���2���1EȠ���22Gt+ �f�3����QC�D[ >.���0���]"�_�w|-�&���I����<�c�̍{����^x��1�a����j��'ڤ�Ѓ����T�ޓ��wRZ���~��dཨICa!Ӽ,�S����L��d+�`7a��F���4���:�I=}z��2}�雳/�6���a��2٢�q��ѤLd��E��G�����NK��(� a�Yd�o3��ڙ+�\��od\z��~�,����i�>^n?��z���"�]=1���A�du0O�\�ә�q�!����K�aڞ�: h�(Ya������X\�&v��#�2���U��o#d�㧖�1u��U}}s��G�`/L��"q�Ar�8;e�FμI���`$ߚ�%��6��v2D���1�Ч՘	������S����'���ģ[�ߌ�sX���vc�����lƃ��%|��X �VD ��=��b3�lt�j@>!���2���ZΨ����a��!wpl��R��,����V�&�Y�ȕT��J�PJ��wl;~��AB�Ѭ��^2j��wn����o��v2�[2E�̭������٧�]Q:����,�adE@�V�7Ě���P>��s	�����2���J�d����d�uU��'��v|hxL�P_�+}�z\y����b�~�㇎���#�Ȃ<H�Ɯ��0��O;�
7rDr���>Y���9��-�TI�*��֨�94��=f��Z�a�X��y1����P�qeB��ڝQ�f��j��F�Q�����b{��/�y������}9KҊ1s������ߕ�;�UW%���`��)��FF�=��~���R���J1���>U��6��b�����0�?A�k!�����܎�g;�	���\^���%�\�@�E�V@��x1yW��ݗ!����iT/�>n�!u�ٍ~C�$E�yk���=�n���HF]QM�t8HA.	(�c^�39��Cl��e$�e4�w��7���U��Bս�Y���Y0�[�<�,uP���_f0�N�Fڨ^�Dk� Pmc�'�We�~��`���^6;.��@RZ�P<�j����'�t�g�a�:bN�SL�b�|��9�`���d������ �����T����S��)yBw�����o��I�� i��Q$�����`�.߿hp?g������Q�Ni����d�S_��{(�q���'ւ�#A*�/b 4��R�[t�&ө�Q���s���[Z�oݵ4�(^h[�sX�í�ⳉ2��1�8y�G���/MWSXz��0S8j�8������ݐ'a�4�Xb[��f��)��D'���q��X�"T����-��g�-�'���W���f���W^P��-bd>�X�1ç��yH���e�L�95k�h.p��}�d��g�H^D�u/M��nŸ)�NO��:��������rۨnU<�h�jcO�]�"� ����j���}���g�x7�ś�'�8����Jh]s~���|g������>gf@с�1h;�L�#��`Tn���qاvy� �<x:�a��C��0��Өs��*�|D�-e-�ǽh�&׎ l�Hԡ�\O�YP_з8+ɘ�.m�����ԥ�KX8]x����RalP��Z���9n�r]���4����]2+��O7����eZ�]�q!On'���BaR{0~	��}cb���"߇�r��U.�0����O�Q����+���3h�)aL�dZ����OX�4��a��>@�-�U��b�PDR;�ƥ���)E��f�GC$��u���Э��n�8��h5#: �op��*���kx�H<�� GJ}�ȇ��j���уA�6Q�V��K�Q#�8�<����	��L�,ٷ[�Қs13ߒz:��*#Ni
����R��s02�h�"-���{�T��wB���Bd�܂�*�*�c��/��j�m<N�d.ES�^1�9�~xa^��u���cfB�S~zԬ�!<������g;��������� xo#E��:ǀ�� �)U���P��Z��K�f7-�B�԰Np��2�(ظ(��c^�w'�d��L���f6,��C%,������Z��Sd��AD�k���8�\��w��9�I���6��k�'��
~A�I��\N�>�6
=��cD~�
�ڝ[�������#�� �-}Fe�ݛ����⮷�BzȮa�J%$/s������ �1h�a�!�r鑹0����ymW�7 8�� Ş���`��ŝ�P��چ��e���H�!���5�F�U!���Ύ�4�(ε�3�fj\ᜥ����O�ı6��'qfFL��ž>[c���iYA�0iEe�Hud�Yi��.�Jڿ�~�̄�K}�E�����}��+n��Lɝ{�$�[[L4�PjJ��a��s��.08jJ�u++w��:U���s�Ơۄ�K�n2�d��"�"Su|��S]��Ķ�F���1m
�\Nf�#�4*XkNh�05;-�JJ��PU�M��(\OJ��|�iLq�e��%v?7w�W���P������{.���X�3�<_�E9��8D��V�[�@'�	?�����s�t�N����b�_jܙ�����{�D����'��G�H�x�]��3b�
�k\.r�N�u[����r#�|��$!Zƙϖ+ �� ���W�.��Q�#�L�VD"`,4Ǝ����0�2����Z���bEg:�o���9�|��k�I�=̠��V\^�1!�$�VP�i�ƞ��d&�ܐ�:A2[����I�:�#[b���f��:����8f��e��Y�%���(��і��/�"�aP��@�c��4=~���Xe.��iD��N��&���n�U{V~����>*7ooMq����-��5l��-�K0}j���(?:Q.���$ߟ�
��}IkNy�6�J%&z�����\~a!a8��g�ߗ0�'�q>��)���J ����1y�UY�?@�w���12�\�W�U�U��i>%��_��A���ڐ�'e�w�
߱?��0�rN���*����T5u3E�P��k�I�ɞ:��i�ݢp֖!��r��d�Ѭ�O䧡�\�HreM�H;j!��L6��(k@4�p��zލS���?�@�[�v	%L��ܠoG'9��2��&;��F9�b��{p:ȪjF��<4��t�[��6x�B�������1Q�G��tC�V*ƼuQK꒓�~��Nh�-"H8�ꞋB|.'Dw�j�Y��6�%�|Z�2DFD�T���="�b^^JȊ������w��D ����#Zu�mؚ9	���1�����z�F�0����j��W;��w�#23�2Q����{1;�6��A����^���\ٝ��Č�������v��m�U��Q�@�����v�J�LQ{�����@pA�=�"wBC��m��]���?�?u�&���8&E��z���j�X��7��k�%O�E��v���K�!�W'M�O4�Yt�ƙ����2^�����M������L��je1r��I=�:��G�vyQ�O���߮�T����E,�qؚ2�i^���ۘ�C�;2�u8sv�����ʋU�g	��2�/vx�[Z2%z  '���u�ԙ���lo�c��2�.)u��mL�hH� �%�/r5~>h��L.|0n�B�5k�ʚZ�-S��^rh4BOL6Ɖj0A$�Т
|�o�"�Lڢ)���"ߜe��}D�S4+}XE� /Fz��A��S.v����p}�$ih����ZX�#p�tWE:.�Q<����C_�(�v���\5]����y4��8J�OiW��FM��s�@D�?���x�#h��3������ȯP�*̜�+��q��7g�Fgk�E;���V�)e}����*�C
�>�8o8n�[1��	��ç���A�(�e�Q:SV>�%R'�K�j[� YLµA�|�ƳA� t��o�g�=��������k�)&�bhg6��2)����=��tͥX)�F��vǩ�o2j�<��P�ZC˓����~��K�a�L�+,�՛-j.ڨ]	6|{�m�$��v��pP~b8V*�3��z~��p��RZ2\����|v�zFd0��,�Yu��-��V@�o��ZՏ�~g��1��)��l-�6�2��{�E.���79��vٝ�*�Ђio�dy�F��O�KK���3C$4������0*��?ߝ�^�)_zf&`�Փ��fl�&�PR }��ّz��q<��(��"�k�f,��Ϧ~4z���--����X�xC�r��(��$���A���!�~�.�J�vg������[���˫�V:������)�[@��M8��ԢY����Dǽ/�A	ׯ'^����1�48�sB},&���XvЁͬ�k����/��.i��d��ʅ���\��6K!���]2!�ew��iưy7�X`���9�u{����޵�viI���O���X̶N�؄CUW��O�mS��6C�zCmЃ���J#��Ã�[%4�k��d[]{~�pC�D�["3��2	!w^?�?��ϛW�8Q�~��ޙ8�w�B$]��Vǹ��nj:z��Ⅾ� ��e/qr��%�#�*1���
�oF_'�K��ZQ��e"\?#v����[Ә�iN��\���}�`���1�t��c���U���NC�zCI��*C�d���F�'Ha��t�R	`t0�����H��1؟0<�/��TT9_7^+.���/�R�����m1V�=��kY�������g�&όPNE0����]�Q�I��[:��:�.�f�V;&Y��0�3�����9�]Dm,�q��Ųh�^��#�lZ�аC����,}���n,ș]2�0�zS�MǍ�Cۇ��fmܾщ8=Og�S%d�`�F�ܘ�����@ǛX�F�����t4���$��F:p␒�L$�������G#<��4��0.�ֆ���=G���W!��Cd2��o��.qv�6��<���J�O$��њy��G��Ͳ�{�O<�q�
�
P������I!�������.+��h��l�y��Υr���UD��>gJ�O��dBn�@`m���+	v����;d671IZZ�$G�i�Q�aMu��Z^]�0��z��iy�ig��oO/��f�/���=\%��ۣ�GG4
V),��-e�U2�g�;�c�,[k��̉�ºt�Ո3�a���"��IM��"��a	���;�u��Ɩs�����5]�2N�L%�؄t6! H�ʰC&c��t�E�?�绖�G�*:����.�a ��z�L��9q�5Egǒ�y_�H��Q�|���Ir0��SN�I�$-�@�` e%�:�M7m��g�S�����&d�������Ta�~��宊C3܍�-���f1!�䯢g�MT��/wxYe���� ��Ǳ���牪�����k��I} 6���Mn
��E��,2=}Ƞ�j���C�Ҭ�H����,�ntk�S���1�ρP)J=Q�.�(��Ќv����O9gqJ'd�n�ȫ��y#�_VYcGx�+�,@J[dg�8y�-����N����m5�i�G�#G5� �/�+<a<��<��Wҋ�Z�@�B
Rz���/Y�'�/@���QC������H�0����nz�D����/b��D3���`6YC=�*���UCQ�N���C���Ys[��}�=U�xS4�8�m�^~�#����^ã�2q��ۀ�1\-��Y�*7�����k���+�HH{c`R��5_��#���Rs`�-Nη��%��*==�d�B��L']���
���5���=5�q�OcN:E��F�.���w�zeO/���/��Ѫ[X��
��]|҆���. �����K���V�+���	ѕ�X�
��6Y���z�
8��������.�k⦿9�2֓��@/�V)��RQ#M3vX��y:�q��5���Ko����݄s}4���atC?Y�%tt�ۨ&}��4!3R�ј�Ċ�*���,Oy��U�$����E�"]��Ӫ���4��N�ʹ�����s�!L�����&��"�C�MS0|nY��K>cc�a�"�'v�2�M��(\��o��eE�z\��#Jt�k[=�4�1s��6��~1@���ZM(D@�ۻ�5��
^�'K��Ħ�+��D�:�u'�����(�T}���v���$�4�g���"�?6�۳�v/<z�*���i�Y��>���\=�}��=i�)
�/F:�a�ن�����k}t��'C$܀,�������dkݕ��NUz��o��Fp'5�?B�\�+Q/�
�b�`"�C����z+׀��$�}�FZ���Geř�=���{
6/!��c��?��!�켊�(�url���<�U�;����OTݗ�C�X5���/'�^�����fdA\�*e�a@����KTƉ��5��w��p��޵�e@�`6d� Ƅv4#���v�W#�*�_��(��D�~T�J�0=�V3B����i���`k�l��3�o��[CE/uҳ��Q�(:t��MArŃ�y�q6{��81ɱ�p7X�������٣���/�.�xJI!y����s@���<���שB��2��	U�\ш3S	T"(b�e4r�cȋK^��6j*S��Q..�����wr�H��eJ1w/>a^��L;ft6������(u����
ž���jǮ�ɁUM�B��f�������I9+�5��;m�	������
3�}��垴�C�N���[��d*��rW�E᷈o�X������=v�x��!
]�<m�rH_j�C$�W����C�ԣ��j|�+�$��u�:\��n�>�V�p�}�
�S!���6nRD?��x��~AuI�+KFT%6�W"
=����»��~����j�m����w���#��(�[2�S��z��O�_<X8��ԝ)b�CC��R�'X���N�%!;M�Y�F��l
�p��L涹z<,��>�O��譿]�ۺE�Gk�U(!R�0����Z�7e��pM��.�"fش�H��0h_2�~���	xO����>�8�x��r��[x>j��ڴ�h�c�R��i�TNt�yY�Bt�'Wf�6�T����<�j<6��Uo�Ǒ3`�F�r�@Ro����\z*;����en�ƌ���X�-o��F�-�>���5E)y���B1���P�������z|ih�����8��Df� �l��!�//���j�2�C�͒y?�hnQc����4k�X�+4A<$��ޘ�}�n����,^�ߥ<y>F�R���svF���i*��9�:�T�3 �*�$��!h!�FЁ�������ȃ�eX��87����ue���Ǵ�2J�w�eW���Wm��զ҇C8�"=�:��RŜ�yA��I��.����+K��������(��y�~��ަ_]q9�	;4np��7�g��2Dӫ�o�Q��q�|{�^���la�[ �$�E�"�e����F��Q�����v�1Y��_�����<L`J�A�Q��DVbh� <
. ��I��5[�C�[� ��[o�����i�������0��q��&��i�]�=߮x~����N7�8_F��/#3c�0t3&�Zt�n�����	��?�������b e�?n`:��Q�I�8�Z�rN�nS%i�~$Md��
��q�g��Rh�������pq�:��=7�ѩ����e�Q3-�Jb��Ta����g@�L�uK���>Y��+�3}�����׸&N�u`S��97-�^����tp=��&I"�f�ʚ.0�����w�IdM�Q����"ÎI�%�N_G���t<����Չ0o��;�.�C!l���x���-�d,w�_��f�߸L�-'6��77�K6$Wp�u����
S�3J D.J����/�h�����(qZA��6�I�uE
h,��`}&khC��S M���I�7�G���ަ��_���.F�{��	�G	���K5��C�w��Q׫��BL��}]ϯ���%�:�y�i�*�`�.�)��P���H�4��N�A��z��į�N��V���cv�%���Զ����cj�O�GZZ/�;�愫�ݟNM���a#�j�	'����>e�xzpM�y�y�����(E~�Yc�U���Z�+	a2 ��	�S�����b�O�(~�3*h���[G$��߀>��r��Į��0��{D�$MC�g�7a���홝���~�������}3Sp�(Ԟ�R�q�13�y8'�1|W=j�=����<F{���Y�c�R"�U~h&A�n�[g$���RZ<��\Q�-=3��Kѓ������p gB�8	���r\i�lm4���Nu�T3syYq,秺��9�_9Y�wa�zh ����C-�4efݷ�ƻ�'��/{܌cE�+/�d��ܮߨ@ma���ٛM�#�a�P�e�(���-4�⧵ܔ�|'%�ssR*a�����?���tH���B�(6�D�ܸ���N���s)�(�{l�	B��y?���i΍j�y��^��i�	,�H�M��$Xi���/��a�0([�W�Y{�3�??�=;��í4�I�^"��c����\�����W�]�V��}�*;�7��u�ޥ�������X�T��ͪS+\>FA�;��iXv�(� �t�.L�}�S�Ԡ?A>=%~���9VE$�ܚm�Ъ�<6����@�I�B_l#s�{	��^�M�i��]"ݎ���O����ː8���	�HW�4N�i>�M�>ly�A�}�C���56�Q�Ox��;K	����r`[>E�5[�_I�>��.b<��{&�k<�'�:GH��W��HyKxy��7V�sH!X	u�ȆuLI n�;Ww#ۈ�k1��we40gz� u+�q�%�d�V�i��H6?D���.pT�q�&u������8�v����Hס%)r��.H ��~�H�7��
6CÚ��#z�ÿ��!}�odM�=���Z1X}�Q�xLZXZ֖�׷���92
i~�G�X�D�.�=��������"�s�#}���k�졊� O�ά!ҴG�>��'�쒢f��8I��l��q�"ŗ8���7~���Ƙs��r5�RL\V+I�m<养*�)-\V�B^����E�pmh�v��JJ�S������� �(��"�g��)UK�����ou�#*��4� L_��Kc��_�8D%��ȭ�J�eS%�G���oP���{*O�Ny����堾F5�����6�VD�;��xמ��{i���z�󰣒&��h�]�b+iY/�^���F��|&��8#*4�YfL��M(%øT���s�s�k�f%�~�e�[�e
��N	��f�-�����.���`W?�\��3:<�&�]��8 4[8��f�8�G��'�֣�9bZ���*���@���"5Z��%$ѣ�e��w޾5�~��r����Nay7hx����-"�e�{��k22�lvnK�o�>*��gg�X��tY#�p���*�͸n��b��Fm���<Y�̻�>7�z��1&p�/6&��Ξ�?��$��������ܑc$�S��r�6c.�(�o�0�Ǉ�#aZ��8c}Q���p�5�1�.2z&�F�@H��.�p�j�3>q�mT�\�����d�%����E�<Ge�U��2:8�}�v&#���]_2-��c?��[5�7�:��vZ�"��ܷ��gO#��0_��^nS2)(3�]C� �)�\��N%]���#�LH����g���D3��l��,;?�<S���L�9�BQ�������7��j���z�<�x�#y��\���-������9�\_VG�qZ����<I�xt���9	���<���b�r�f"��t��I��]�� #� �1�MC�,������p��(���m5�M�[��*��+���gHj��_����,���Ϛt���Ei�O�ٶ+����R��g*�F�+U���F��Wg&F�K�YPPM�S�sp�5(B�FO�@{̘�Fn�^�Č���-7���|~��6b,h ��֢�x��7G���5��d%�E���B�2�G���{;RUN��Ե���p�V��G�,��ϣ/N�!�Ii8qE����Mj�1�㥏��ŕ)������*���L.Xb��8�;CLLQ���)_#����ߖ}��~��q����z�9?�����O㠔��O@f
N�{y����o��4!�/��qy�aa\�z�fo�'}�Zf$c���K�z����zB�hJ��}��᳚c�_��2Nϛ����,5�vh�h,5	X],��Ʉ�pz����2�V���μO&UO�!��C�چy]��I:k"��2�X�_��v�f&�ph�e'
����~_MW�n��n���&�yZ�=�5��@�)����:�+��N���iA�,�נD|>s�tĭ3	m�w� ��
��V�<jB�x+�v|�T�l�^���J�iN[�����`|L�ĩt�_@���I7T�xoP���~7m�f��_mW�2Bf�]�� �
{���\Y.�[/
����@����e�"���m��4�EI���Q.5&s;�G��<)�10=VS_�Ŀ����w��U����d�>���&U�R�K�˽�������>Խ�H�R�A��ߒ�x�.bx�bt���b�k*U��vx9�l�7U�����IR/*��}K5�Nv.��+�u*���q�����Y`���U��Ǳ�����/�V�
e؄���Q/!��V��P^�r�¢#���O��:��EL��(qS��T�0�lk@�jQ_s�g��)�fvr�-bI��m�	�`�_��.���M~=?���#4��-J��V��1��Uf��5���y&�ͤd�5���/c�<3����<w �͙!���zB�8J���g�S�۶��E��W�S�2;�_�o�,���!B���Ͱ���Ȓ�@#΄�\\�ǓF,v�jB���\��z�,��V����-�����)ۚU:\O9�R���'|��l"�\�iz�g[_n�c�M�w&�T���F4�Yl\�e���3�D_����CK k�U3�)-2��4����k��`!Od=��>*&%�kPD�~��T�k��#��t��i(b�μN��~�ӡ�������8r��ӬE��C�ŤM�ڮ���y��+U^���E�B��;�:���!�J� =��u�͗z���|��7��ևR�(� ���we��e�����R��җ��UNۄo9��%`�qDE�TJ~˿;}Q7i ���[7�`�9A��;�nfP�5Q��X�7��\èj�t�׊��	�{�Y��>�z��BM!|��O���Z)*��z�0�t�8��}��j�ZLҚz��ҢV�������i���`�ށ=f�f1����=G�����ǅ&��*�r��%��;H'hI�/0�Ŏ� �t��P H8�J?9q�����q���� �C�N��ܶ��l�c�����"�2P���*����:��g��g�d�o;7=kk�*�Q{��>�_mC�
�Q�+Y�ń
r��܇�����Sߟ1:�$�����!磚*5X���#lg��
�m��:j�.�uHP�wĜ�W~[P��f"(����b{	����"
��������/Q��:��v��l��j=(����{����ܕ���Z��`�,;M��J�mV���c�7P&/��Z��R����P�T������W�ЭI��������k������(鐖����j@�r*��x�jCM,4��N=��M��M)�����ǎ�K$r�^S'I����X��CG�?{*u'��3y��v��L��sʸ��3�ۚ(��rÃ ���ؒ�L�N�Ȉ/�>>�A�]BK�x��	�����JlP��	�]��� ��p���J!�Bj��2�}>��B�k����>�g��`�k�F�b���\K(�Y(���6�3TI����G��&ؾ�o�����Tv醀i0+����E_a���m�߯�OR�/^|��0K��*� [Dn��P����v�J�u���0��'"�D�q:�6m�&[/"W�j/���4}�s�Q�bV�����^�2�?��<i2���Ɩ�����w�˜�ŉnr0Ȣ�pTI�.�]ORW��e�2D�5':eC7��d���0D%���|@PO�
az%��Í���[c�=m��:��#D?t
��Zm��P	�˨o���*���uu1�/��f(�Jre�>�[V�GX���F�6�� �Rl��2$܊��e[2����W�htb�ih��íJ}�x�Mg�0��a5�{G��BO��e��߳�f����M��K�����-❸k���[ћ�XD3�	C�s��F��B�;.�<I	HW?�_���v��,��C���rH���@�"���6�ČN��d�h�G��U��T؝���*u�B�wZ���bK��xN���u{m�S�MɊG������Xdw�˭�� P�>���J�٬k>����Y��D$k5H�1�6lm�ǽ.�&�-�wg�Rr���WJ�Q��ڶ���I�n���FM�I�R�BI�S�zQ�Gt,lhң�o�[(�q�9�@��	8:�ͪ��US���ȇ��$�K,�
㟩q7����7���K���D��fC�PI�����.^Y�%�4p��{�z .�{��VzKU�D;��Z9'�3�����Aa�5A��M�S!�����z׎3�#-�,+X�wk�,|�����92:�7�C�	��o�d��H�NB�_H���ǃ[M(��ò�d�.T[��ӕ�� �+�#6h'������ޏ�Φe��(�_-�P��ّ�N��`^���t�s�%ׄ��<Y���!T7~2m���݉�c%�t�z��ׯcԄ����@�K�F�${I�O}��ό��t�<G�8�5GUd�y�;�Bh���d���mj��`�30I����䓣b��)�Hឭȝ\*T��ϣ�þr<�N!�z}�1�Gfd;N3��;���y�����R��KOu/g��>} �oQq}�l��1���_�-�bx�*^�5�E	�d��+}���JIި�OG[�3Yv�}�w��� �8sAl1��yc�Y� �[�j�9
��ä�`
�!��;h,)mO	M��m/Jw��u1U�u_?�*��ab�R�)�Ƌ+k΁�����\'��4$dx ���y'��^c<�y
co�)Ȕ}_xbk��s!���9x�q�ͩ���v�@��z���|-�1�"����[0bx5J�����>P���ݧ@��T��u�Ӏ�`�b��k��)]��ꋋ��iƘ�`�t�vH�0�)}}��[m����ƶB5d����}{z�H�������v�<k��ؐ�^L���> Q]��Bd�s�?8_~*�1���Ex�n0<���ލ��]�+�a:��	ZAt���=ZΪf�����}ZK�0�(}a���WGh�k��5yY̯�O1��A��4������H�m)�}�j	I�� �>���ɪ�N�4��*�J�/yRE�FX�a>�y�]�FP7�И����$�p���,��.�bCk�����㽀o�/w�)���nҋm�c\A��a��1����Q{'�A�?�n�ٚ�3��*�f�_m��;�ңq�}Wx
�N����'�T��q�r����u��fg��|���km(4�AP�r�'iB3�K#��>��Gw~;I�nǻC�]�V ���D�-�+��*o�1=
te��Q������F?·G߽��Ιה�1ݴ����P���#����t�3�[9�L-E�~'ga
�ݳQjפH���QV&��o��������`F��(��t��zܧc@,��o��bd�X��Y?9;Q�9�����~��\�K3'c�D4cH�>�����T���~O��6�C]��xQV���7 9��R7�:Ք�o��X�Ʉ|�9D�Eڤ��,0�xLOb�H�L�<���W��; �9cH�e���lfT�]j8s�������jV�J�e=� �3F&�����'��)|��)�`��G�M���L��,�9�=!͌�����(Q+�'E� l"Čl�,���]�7�tǁ&�sh6oFT`&-Jvߜb_����g�������ET�%�^�S�.�2����}�����%	Xc#�@�
{фb�S���q��S !H�9D0%���wv�6�|d�>�u$S����qH�k��EE)َo�^S��8}���҃�fk�_2}�ݰEoey'K�����'Д�,E�Q�X-�=�pe���5N��LFsbɣÿ����*��&R��_5�@�yb����5�伆��K�\y����|�W�\0�n��W�6��������Iz���;�q�&�]��AA�����vTQ����G��|�}X��AIx��Ž�a6�ǌ(���C�S����k� �i�$q�Y���e��-uc'j*6���a�@��/b��f�E�u�����H��F��F���\�C����ˮ�����4rm�?�eHK]��M-��� ��C������?�/�Җ���&ԭ������ܭF�����(���L�|�J�Q��,��.M_1���B�^��ݟ��Z��� ��)�c��c��QWX
$o8��.�$�Ku�'Xg��Lw��+� �:�>qHm�<]C�PT�&�/�9x"��#����t�E·�z$f���f�K se���"B�0�EaC=���H��O�q�#V8�
��H�ql�W�%p�C��Mݘ��$>X�C��̕m�q��cs�>�S�\�d��?<�PF������