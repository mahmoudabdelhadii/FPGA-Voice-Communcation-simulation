-- (C) 2001-2016 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
TDBrZzGIKlc1UDiCvkZSqm43+5rvVsjqsuzrvtp6BDvzZiWTdIMSbOTbvwXpRpt7qIk0V3JDen0R
ZMyfke8H8BhFxXPiOO0WfmnbJnMBT4Lp5sdX75iqaXTOWd7NDthgUsqf57ABuxkzhARav//nDC0U
/63V2rGLem6AlJZ0g6k/HoaqwYYh2GRQgvRiLKCkX6lXqkeJudJ1r0odkil3IN9Dis0u20jjQsRh
4zHJ/ZUQSrsbF5sxesyZV38L00Ss8s4Z0SUdW7U1MH++v/iVo4mVWRydHYMsS6FvjqthxWzvfhGT
4WmU+whLPWfEvEFu36gA5piwJgH7nhKlkCsssg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 2368)
`protect data_block
XNPmhmi7xrvtP7VlSJBW+4iqnk2nULO7IjAXL1qsgleCxXKhFzLhhEaGp+qZvzXEwtGJ4qRV8XAV
o26awjaKriF8MZerQF1Q27qpENMYDT0Yp9Pl2pAuDpfm3uG5NMmoubFKqh9bZT1QM3141G+PleXr
xMZQwjgh9Ji2MebEqKbBCfON2ygmh/sriTMejDcpiPxFBMwYgUO65WFWGlNgu0XSaXj6KGSfzpDA
nYTw/DotfG7p8nEhBpRs8jI7eWX9eZK5/AZ4/C4Kw0fBpTGrBIe7TpzGfTa8N/EHbTAFtxlA95gA
Qwrmff3est9Ygr//7Zg4NM3zWGBiFe5SMF5Euyfrxps9tLXO5uGwhfJg4DaNLQP3p4vSuDw+K12d
atLgo6HvkGT25+jxU2j8zOv6ndmrChqIxOZun1F/3KRj/sn64HmLLUPST4f5RkQfRFPX25UVxw9n
JCUtSedTe25hTsiTNhDFdNQJl6RZ3+RU95nAPdn7C8czXMuc9ju8w7EFrHHuqHjRoCIQ1Z5CciTp
oE2wSVVybzCdkXxhM5a1nyIQoYkdAINaY2IRefcbrJqDJbQYMkflT3XVz3izuSwpI8iIdztvf0eo
tBwAqHR82OwdRsnUmj2exZWO1XyxH00mSBc9BPyzwiMEGfrfLP+H3X+mFxhTxjzLlXHDKZPYBnEb
UZYcg8js0ptbseuzwMpfAhZLNsFf+XBVFM5i5WGoJRXb2CPSH0BHeOTGTctI/Z1JIFho9SI1pO/m
J8pLSQ6nd17F7e0Epbh2b8kzPqxs65+l0+Wcog9S10hjZ2dfJ70d44kYpDWRzaD2pn6dKUqpgokn
tiAgSBqqbGiZsk1MlhdzrZtmLtnVUL5iT9byRzDovCVoPxJzxvz4hgqQbUGAS5eSRmIuQ/P9KAYq
0zlzlsji3sX7uYccayx4/ZHYcDoRJRZ5L5M2RhSEGZ+j6OB1oPyDkPXbpiV0fYmbRyi2XZwo+lLt
Cs4rcW72paXZs7/0aYkcVYG+wu7wsjHdz0fvf1HHeKm+Moe7TB7aLSrQDL4sIBpVhtuGpCWWtZXr
PvJSzV2f2Jebo5YWGIskcExsrtvh74VC3zsanc2sUEMX5FGUsSHgbGtI0Xr+ZuY+3hb43UevUNMw
s6QkqpE1l1AHNzBQVar0QUzqumhtEz+ciJQiaMv7Ce/RmqRdYDEBxILXlGkDAhY/XHJoX77VuSfm
426LGbkwjsqFg6PnFP0EjbwvXkzSGSxXCjNOIvSWeFTq7//jpB1P/5EcNJhn/u+DceCgCjs7dUeb
4QYNz7dDX8uDBdPKL6leI0Zo7H7Yxp8gjsfWwKIbpXrQvhhNge02Uw7P5CWQErxerGDWGgcvpxT+
x5R8T0xVDSd0cVuqGQXhBWTEImEYLmg6pA14Uxjtyjs+d3J2GlRQtQmKA7Q5wNLPgOpJRTViqoo9
IGCKy/v01KqjHkfaCy9KApKwVt7JI9fdbecb0pBAaCF+9RaGOjPbEtA57DytDw8Dq9sVwQhdlq92
UBqdgShEoY6PeXCYcD0sNAd/HHJ+N9OrQZRMxI3hCpM0nOTTWtArsO4kOuNl7qsCbogNp9K1hXSg
Ci1Vq9Haw2oi+EOjldU+BzuC+0bUj76ouHGoSuhM+oOvU5+mEaLdBJjmxf6edXgwfiwT10czBeXR
Wzz4AEQSAZ5GOIlrgohPoDDfXe9XF7+VG0bAC5qeoiaYnEdQaMBn03L09lA2Jv1+rtONVjutKdEv
XnS0zOudcQTU2hQZZJ+ARI22Xmmn+6ZM3P1FhiSIhe7Cc0mvjwYBMve+CeCUjMVJrrKCCA+c6+SF
p8fhrREXZ3YnbZmdDbzyF20ti854jTFLU/y3nMb1YCkGMvkVRHX172RFzUX8bTLAIXTjT0sZxAlM
u5aohCUyg6tOD43y6AHZ72ZpFkMrgGR/f4YosdUq9Hk2PRDmU6JcfuKD3u3HHDuaqkrhOFdeNyJo
LjvaUfYYY6FHLyV0KTLWBbQHWxm0RH5DZ58m3DZ4nfpD8UiSy8zSDa6sOvfpQEJUofBKcLa4kPo7
kYm9KxXWEo/5ub/dlM+BMtNxPFFFJGGwHuagLCGQUcMO8Lun+UyYB+rGqMttpprP9FM3WULPctkH
rR8LNJ1EuJaIVYUJzeGcN/oXp5Jf59jtmKMbkUfcdf11bfujhg/x4yugw5I2VMiStTedT/1AIdLR
AZt+U/98rqxjTfnoM089PTCR4bgR815atirexrEPyeulv6W+2CgPq/2DT4Yg8veSgJ07kmz0FI+S
6nFofwYZ3WfeG5833KaL+W0tM/tMwqWftv+ciIxfQd6cd6Nw1P5tsbv3i+qhJjehqsHqY20ZtIUF
/coeOLIF56QN+kpWrECG96KEY5DgwMd6THEQh20ULPqqUKt4HZeudc5GKPh0kzdSpzq7GmgI3Txj
jqHX0scaGkJa/6M1P9vJD245OO2M2K4jgZ0ZWfIaXOJDpHzvbdw4763+wpwDpvaUPTrZYywQDnwg
I0InrVYX4hnvhtWTiRBpjNATqYLiRykFdCLMbtMe2tfmnvvKlhGO6NRzEajD94oGOHHgKxvB4E9B
ZuAjBW93Wkv7YGMwWbWlRMwE8Xw+0nZ34gaL+1wMEnKlBx9ZGFaf5SP/YnjABlI7zfMggBF4k+us
gfDtXy7Ek9GTDFthjKygM5ntLIGByHy8YYadGY8eI0ozq3gmnisZH2gQrOy19+ZLoAmOhAEUfYae
bmQkXix/xd9A8bHG8dWGWr5ilu5wRoseVLyghEjEDQl5kfqaCWletc51SyqJAV7t+wnpUXB7wDjN
oDzSA13bIO2vs8OgamFd0cPUMG5E3xDaNHCQTwBFmuRxHfXSzb/KTeQ4RfXKlWVZGWyZL0/ObLGq
Qx8KwYbUBNdgMY68QBE/ajwFc5cHieFyVPbfe7qpqDfUfm7NLzfyeuRYzy81QjiRt5PJK1/GueD2
dwFZE6omcyTt0rw3APlTio9J2fgYva92kmJwUU0HpsJR5pLPkS6g6sY/kKIxe2vG0cbXcP3al6BW
i9vKMzrR8AfVgippaHbwj+N/mgGIOEsVwfkVi78CVNmCoavbNAYvzz3en15ij6E/9jDJnhHhxXDZ
GKfPZxl9yYxCTgolkKrrM1jgsNAkiYE54ntcfjo4kw==
`protect end_protected
