-- (C) 2001-2016 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
SssOrSCckQKEi/Q+iirVBZnlGzzV810AP8Y1++HGJAnqHDvEhcZ0XgbhJVCdaCFHXsMOyiJBuheL
6fGT/GCMWvqwvA7cVlmELDheqtZckhDH6wsIGFewIWhC/m3n5PHv3NlAhhuLetAQyIECkglqpNkl
5okiqS8FvaqMtPBH1/gfm6jdSYbCbX+YHLFupNcLBEIBhCF7gorpo5wmLaVMvGDv5epBwnS1rcM3
64fWxWZhUki5x+/1A5OxYM5YNpHFklsAW0rSATZUTlMh6jCXpHE571djng6Kh4dZWp4RBXnb1VZZ
/+uqgE+bCPMmHKmcysHhhc3Zte2eegW8YwAdcw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 11616)
`protect data_block
/988DVzBcu3mQX99mkiV/+J+Tc1jVDj1l/UuFsscrEXw7/XW3X/IXHcyxk798nBGHeHhldPDGiEL
WT4F+yoUtW2Y+dOjb/lt7djcgHX8giR76ZPqjKBUVUVi+8k0hzphDp+T7+oY3xPE9JYC0gg5lsIH
boSVJk95MPm/h67YwJ7aBqeN2CqxIyklvq2cR5eZXr5oTu1g7yOyc1n3MuMDgrxcgUJVztaNbQuA
ZW9R53VloWcmR8GDuXj0nBU3FyRu4LmK71ECH3vj1ducQhJX5cx00dAwayK3BReWHKMOendKaMHL
P0qzMHKfpuBHO90WGDUklV6zyfBKsORVdasOKydENNJVh9OC/Wtj7ep0ETtstdiZyT5n231o2aVF
TEXM2x+EgdZIxweQcJfJyxlnSAvxG5JlLTh+edeEVV3zO0MLVodYouYsFXZbQYcp6ANRcJq/g55y
sXmudrW6wg9OZ4uMBv5JuNWUbpm3t7nYylW1oPSqrYmUK/tnV+TdPbi5Fv8l8scgUFSbR0Xqt9Ng
lvOynE0KYxN1s1Wdq03ZzgvKuRBUOrn/c5kjYiNNZnUDj9Sl+Cj0E/O8s8rYGMwIIZxXPogVCteM
r8I1YSZVZb9vv1od2/IfQwkUW37IAlUP5HErfBWFuHGRf175ouhagRQ8eS+H/zfiITuRGPnGn5px
dn4JHvjd4xrpBMZZ4r57wAUmCEHqYmHfRzYfiQeRjp4mK1U1LM4xnLxEz25ac42Dp5xlQji2GsGm
t23y5Lz3I5ORkmWzOzaAoIh0P/1jVLhj1V0iPDeUMxyH7zppFeAkRW9WBfeHgh30w/tPmp2an8sL
38Nc1LZS2TqN9aUujIPwK+U19mc2DxHYCGgkjzEzUKbijBflApMUaumQNY/sqLvoOPVVXpNdSzgO
m5NjR+geP5wW9+H8azOQsyHc/uBOb4nMvH7vLHmKtb8SbmaNQSls34ubJhwOWLFCFasoyRggAsxh
6IjXcs9ROdwll60lXXoADx6A/yD3snOLU3YdRu9iNKUYWEsSZUDMf3Bp94JO0JbxEzx9O3lY8LcG
Ynfik7m5l57/4kwgsSBmAKtCaCAqezMs7CGiTv9QhzAFC6siI7yBPkr7hKDZoG/ioFfoPalajYt6
inxZacFa17nD29jsfjWaeCQ5w2Lz93u8seF9srbEmHGuGxAsgVk25EMecZ48xBe+nQLDlslkN8I/
WBSHcJrSWsg3rsTKYT6KLNnvAoInP0G96PsE9Jzwa/EOnH8KydKWJY4TeNmFa5UCe9B/yy1qgnTm
6JpeGW45xVrdcUHilD2a5YZGh6Jjr/bybrbWaBXGEYaCYBYqPdPuetJb+LxoCKbQbhVJ2+A0vH9Y
TEQ60KwdS+dm4hOSJuKx0R3PZ3dvrz/rARD8DyqCO5nmjrhH9AmQedPO/XTgdNyfn1QGXGEBes9M
i7TgLblbHSO0XrRFZUzmFVmE8QEziuBTpxp6NDFalsBurYLYbhE5oSgEktWLOE+ElSWQL8pzjqhM
WZj07fnJAvjWHDtXekqFXXtxPBdIrtTHvFNtdcb8b2n6HL54h30Fr0Ko5cs+u40nRGb/IvXk1HLw
PsMrmcUCp4kbtRHfOuDlh81k3JmdUSQs0wP/ajDLa8fgqDHVnZkB7SqhfZpv+u8vmM3glORga66C
reo8iTSn4SyCzEHhbQ+6QdKSRGVkAk7nxqwjrO1UYN3syGf1s9TvptOYu+UI9rOzAnHeRH66s7qT
+PTdQeAhOpm/BAohUSOJ5TS9WDXjkgsNXocB9O1HPTbi2taM/7/h9UJqrG4RO418VH73g7G1cNPO
JUgxaYhO9QKTJhIFaCYrFjGpZGmM5WbKPxGaHgf28jYxJtJdaukwLrOW8E8Jpb8xVFvLy5eFPBZI
u807hHvSklH4a52zZNpb6dDHEwhvNyA6jUe7P1l8+XmC1+s7rH37rZnyezdDW8c7ASUPGPpXroec
A6iYMjkNEr53ayWCfpg1sph9JxbPeEwMl0wVpRNQH3mcas2uu2eitNOllG1oyYFLNzO96Zn2H5qS
y46pSz5ebD5CxcldcJqKA6D6JF2kh/2v4NiGBMaOMARTYbXCLXhoUhWQdNB3GzcPx5UofxBh61Dk
8NJPSjQMWVOFOTOZSAv46L5RDjF+LfMA1IRX2ZY/sVtMH1HCSv2MlpT4j0dS0wk66777ysc/aiIF
LtidB6mcT/d8BxPPyokAmQY3XM+hGZI8nzLe1VQorpkod6Ya8cxzw27jbRzR4+CoL8b/K2y2nDNK
lGKPiVSRa75nCjKMg9yCv37EbNq4WDimvTqwrTYkUdHCJ7UWDuDJ5SmPknHR6dsfz2kHuqAcGyNU
UKPSqcee2SVT8orE3YIT5b5ehQHUbJ2YiJLTGTD5LJ5703upGXhHIeeftK9OrHGcFz3TNlw8PMXZ
lhKYZ143ySjvxU/3UFUMtIQiQ9pvNP4UdhxTfH4nWh9CdNM2Tgj/i6bOK+SyNoK6LdggjC3IO4KE
bl5g5MkXfoRUQDEUGIjWFKPkQf4M1WlE735F9Ak2ZvwkRd8pKC1wWxm13nBOtuxxGC+sXjiU7skf
sNJ1h/Wsb0QgbTupHvTaSBQtRlqeSTKLeaTdC1jJK+NnLsMj7m0Pj2DzJa0/rkpyC42qvS4jWzo1
UGgsV6/Q3WxkiCJz7XVUUkJyrKtydjz1lzHIkGmZHNZOzrwTAmFzAKM1h2JffLw0P9CelTnUVb2F
p3Po1LZU6jAU1LBb669zBvp/E4hj+y7f5FgFBzratWJc1ZKaKQEOgYhpUMwc91FRfa84s+mTw50V
KAiReaQivj/56UpcgfusnX+vF16hLDf9OuCa9NTOWgqvQxnsmHsyDAZpWsm8LtwbhpW84qoGdy9Q
yatFOYmuTuyJWZQhfvvi2I6owhccySCeCOIaDpATibBne4lOjeyB0MTHzUhfZCs5PPVR2G55W8Bw
1kFzbfWTKtUpP1YojewSUnnHwScfuQXMvlDR9Hro0WsCGMXBC1WY2qr7SeUXqAITbNwMJ1NvHfza
3VvcwlA6BDr12no0ENZpNDAdTcTHDGdb9IlBU/l/J2I7F+v8UN3E0k9rHyLen1foyT6jHjUNv1ZI
PJGrsvV2R/EL2tcl9ZFOndNtf8lsuMHR+7f8Xs4/1IbGJbvU1y8UmdWtDuJGzFR1d00yW57P2Q1H
7ziS90Z6ePorXcyB4f5SWZuClPdKWILC+MZDaREEGzjULI9rd/dUL2TunG3nhU6Gr/vGVevNxHhG
Jz0S4JOwb+FmV20WGYTsdfVsStRcQ512iHtyPZ9hoELr7NX+nabMhZcYUelJ1Jjoz9DOe9zHIoib
uczyeh7ozSIRsIydQ6Mv0rK+CiIUEmBi9lexWb3qf3MD2QATXQaF6Ixyf/XTLuiFcXFLKXleLo5g
RvbdJMdbr8VQQfEF010c5ofGoshEZNCo00cWFhYYJgqcOVA9qslWZZPvL0cFc3bHkIeIEi6k9hn5
lBexswDBk7e6GErvROVhL4gnkZnBK36pOQivjEI33cW8ZoM8SWdLxqmVb6siOkUfUKWnGPx2J/Zw
qP0C3TgyG13RNwE+YjblwSMaraBgsBZsPmWcwe2p3lTM4zI1MzFxLuXrU4xP9CyFu7MI3F7msqgr
t8fyNUH6qkZrN47gXqQdyvWkq6YBirMEDnWE3SZqNRkiIJPDWdniSIFe7K+wds/LFzGlDUa1DUXu
UMnJS1irbdjE+LObAENh2QHyZo7EcIqbB/WGRYWpnrSeP82tWpfG29uk0W0fzvcMz3Vstk1YWdsR
c/+FzuSYgJKJUL63iqIIJTskMSWjrEy3dtigqTEhw4qQDSzagjCcX9NTvE7fFQ/gnq+al51yGzjy
q5L8N7E7yjhC8JHcWMAo9EJPcbPUSLAAHMCvSYSB6pQ7MwLJ1AIKiik3V3RZhReaoomIEXGIZGD9
Xu/z7zlee1WvHIFVB85jqJQx5kyVfvyPUX5YI/NFuLNFYS6DOLs8WIOeE8nJcgRKo+pPcZjvAuPj
2mWS5TDBGQA05nsNeiwh1llRUBVDiuHFDFBgcPCZ93f23aNE0swnqQ/OH5eNCZXq4CvXNgky2Ebs
WLIz0PcCFzSAljAOAOZNaRG0ZmNP9JvLrGKXfrO0gVOoMlon5FwUZAkuVKeln7bFuPjYjX1n3/DE
A18ipGYW1a0MOJT//9JLoPFMP40DHPXPQbT979omV2pZ7yGu7QEcPavVcCXe9hTeXdCVSDZVt9cK
BeWd7KeZ9DHB9/RhpO0oOjQ+BtuUy79mXsSG6K80xawMRTD6jHHp+PgL9FTiqtQUdb6Wg/i/DqpF
DFdUn2VF2ortNRuEVpqpSPu6yrSUv24TEbV1TgcxPzvSIXbd5vAGcYJaufBYtNMDwgJxpiVPZMgn
PSClhELxXz7SF2Nhx1boSh0j0PXc6I0HgAAv8TMYUAeiT1bzxCpCxR3E0RYqI4lRHktXVvK9W4/5
R98fJwZuQ6oobIjxUWp4NYyAx589z2QU3ZQG+BWFSgS07AydSJG/Q8dX7KtHWhJ6ak3zGik+wlme
I9TRwgxe/pwhcKFBE/DAqIEoTfarTGcnaKzIzF8esOaKn2v/rJKjjv2X1fXxrsvw5HtdnwchPpOK
os4N9yYHlfdwQ65HVEWB9QFHbMM76038wbnDb2H6FAxgJQpva9lkF48JsFQbP/wu1Huh/uh1qW1C
bwc13FDewZKwOrwF5/f3iBoxm6wXGQX8Gk6oNJnZ+y+kCCOV/B/Nb6l7pkyTV8SGiyhs5k7RzfrI
4qSQJPRJD+SQZTp26rM1dNEPiTi0UYO8GxE3akCkX8WWnoRCbetoMfgk363582OxoccXqeFE/Da1
sqhBiN3gsiqkzMjC+mBBoL4KcyVhkJ1B+T9TB1/HIUxpfH79fFQv4/xOD5tHktVU5Ip1Pka9vo4f
0rT77Q30/5YJRHOCk6kfT5t4ad7H27kbAuE5pT/1JnvQR3rmr3z+a6RksfapDAUY12TI3qrYe4sI
EHUux8a5n/upcHwHvedaGVskHBy6i05BgzZFJVWTJxMtNFAPLncjKhJ3CTXhZR7lNRZ92cqCKeI4
MUGGF/7F5OSFXyW97XaOi1ZizHiXBpA0WD8xYaUJLoJQ3S0/nNPjPrx/APh83ThHi6pZ+v8fdwNF
qS8JphsYJrWqMIqdR2ddBAK7wE++FbTUGb0Ue1JUFYCox+pEYDy7Xea8+9lG86Ql2mxWNi+BCnrg
GYqUGAKvnS/mtGRfJTbaj3TCTzzbmZJqxCRQn6VRwqaq+WR22Wm3v53Ti5ffGrxCgNHmV1wV+bF9
ZrKjzsKY1AhgIrS9GL+YjbZZL8n21mywkgM/iM6Y5DA2gkduU/1GzRxB48qwl5jytm8M9KFq30Sk
bptbVp3I0oldLp4J9yBWZ+C1RMsrjrenHObyKkYx4JvprznBrBIC0TT6r0/mIn80d514sbcXzyRf
7inqeAyt2GSaALFtSYM5s5j5drZTCjFGauLcV9zjEdwf1HHs4ShEeNe0nbalORvVn8L/9+bcomwk
PiVng4gLifM1nG1mkloEtEIWihZ98FLsAPWEau6a/+wL/xBBLRG/ijyeTz2Mrczjf6T6tnQP7ozb
kbLxCmKI3YWDU3LRyFYaWYBH+XOaor1UHt/u3NZG38N8OmPyb6+dYDbcb1kEgHelX43oVqIMDMw6
iYQfWhxHJcaAkqW3Y6xX8zqzC6Vqwszx6RO87mt7iBZPDceqiZrXoK636eFJklbbk7gOujVVPdWK
f/YDbuY7A7YSAWPl0HFoWDjuUphUDX2TiLsJDg7czUSPifKHOazfpJlJpjv/2DYS6lkZc7e+3WMw
EMAqoMupk2YAEMtWt5Tuk1csUra9EivRrjeda+7blLWp8NUFIoL5BudWN6DQHBmaeHEfGAVhlOHk
QKrt3tEku5WPWRhbsNCwpr8KIil0utIb0XKy4fV7KXtaWZortqBWNSuQ4bgwjZf/j4jtyL6JJ2LK
I+vTvpPu0l1E2/6PwRWw53GalfuqwKtC0C4aeHck6jlOL7q4pcNF/kjqAe8H0eC96e+vyLYOwyS3
/xjmh5UHPwTURn39WsBqGHTMGAvsTnoncPfAlvwxzVm4AVtt0evaBicKP/rQYTAl9SsUilPYt8Qo
mQR4BaHPHpvaxK8NxEGeoBSOsk6HkNY5ZD8YajGpuOQRyDG6ZSBxxv521TThRZj0BcYNOsanqKyY
LiCwfN/4EaMqdwbPTKkE7Bvr3dm1BaFWij4/KAIJX8TCBtAlSnavLtofv1hjjQvUbi8c1FeAC5OQ
qN5PqLgdjk3XCHzDGYgYadVc71n9rQs8aiWJTWvMYW2LtIeaP5dyr6La0bnyFPOsJ4s0/NBno0oq
XL+SwweZ25wgeb/8dTQWOClODL/Xm/CahQBamdWNRUdJvFjN8eKzi1vJ7jTGZTDA7oDXHlj6HQbB
JYQUeIFL2EQIye+hDqjKP2si6GL7J58ONvueWqRHkLfCGBhMMmerPUWBynqspPurMNpgsENK3B6T
6TZraNBJ/95udmbSHIHb6IFQZNM06eYHtB0UY3x7wVbvvxHko1TUvdq9dWwXKnBdXW14WEqoGCZY
ZyT9W/INf95Rsr1N7lubYw405tmg1I93boPEx0jbi3yxlurLjIDbW49KumN5ZDkKs2YGfg/ROpKj
J8/Qg6p7jKcs+r8lUYgnpZWzuVZcUCQR/AFn6l5+oPBe98W1cY0ul0VkxlHKiw3cwiTaVc3W/oPc
2lXC3jVf/93B9dIAoElVFXAcvVAM0gemqCv3dU5UXa88er4mBwOWLilsglnDWyvLM5PJpJYzZ3gZ
g+XVN1bJ2mffQnC5D+6SZJrRsTtWTyyKHjJrslanKbFLcRo2Eaf9l4wXRxRzVjr3qtpquFe9Mo3Q
2LVQ1kHhGeWHgk8dACZ0yUQpVB7hjZ+9xrLb8C+DnuaZuXwyR9Ui4xsrPjz18doAZFImDHyXCoYf
ffS5bNJFM/cV4syqR8rTXSFA5d/foOuX7fKXLyxVK4/LT3Uhr9AffitRRKLJ1OT0SyAZvo5Vph+E
I4QrYEf6t7NyJRAEZcI5VyiY7zeIWqXke8cIE48KozQZyOMt67JgeByjzo7gI+UoCw4FRkC+p8cS
RG3FVJIn3G9e472rKl1cZPYkWZmDrea3Qmg83diYVjruYeRwZTCB7LpdaA/Afmh6Gt/Wxu4d1Kpe
o9CeCyxXfljE75D127zG5Jb8429CTkOAwtqEG6Ozsl6ufdJCJjsS414hM6ZE6BTky79jQlkpKOfV
DAoPht/KkNiSDlbk3MBsdw2LvoG4NZB4zMV2W7uwnPbVsNrpCZ8WlKDyhvu/Q/2QeMhS/nUey4fn
MGjhuKr2H4mJl0TxUU1/e/Lrhg3nrnWAyLl36E3+rbRBPw8CBYUf+45V/6XM1ALAzJcVdK6e9Tr/
+1l3Xta4yzA46VzkccQY0jEhZNQxwRJE3+jMOE/H3KRweB3doLyKcs6KWRjCspUg0JRt1TBJCURa
YZd0s/+Fr4PxyZ02v2E/WW7qVptxWSorjPIziQ0jMNw8kCNR1pnNxo9iZqNKbn8GfYv8mLx/KMRr
43Q9J06FopVl43nVUIq8hWcTCtb50k+WufyzVr22c7E25BPpikky5GyCjHaSNrmbMM8PKa3+QSIO
oNiNDQhoG7VmVYWCwtyvs+f8WLbOtz0WyQoWlQOiU9BMtj1ip1F8IaBGkuTvgKn4LI4U/msK9RTO
Kju9qrLVFMHZMJM27KCYYYRUZY2IJRCeVn/1GiulZgeQiWTZkZvAiN5JjWh4a5l2wGxcQMnDU30I
Ql4h4zh8iTjhN9QU1Lyf8geoaFGPET+uHp9o24TM4X4D5lgAQxwa/zEi3WClPVfBS/YUXdD12yvw
82YC2P5Fl1VoBBo12O3Gay92BTL1mHYchuhF77ZCzIzcH0ATlXVIV87PawnpcazT+U7GSWPKLoup
IyQWDu+xmW4LqdgiCtWxaF3jGl/OfR2ix9aOYBHKjuCOhim+dJFjdtCw5oI7lOZASQXyR1eRplKI
9dKQEm3oU5vURUIVRnXw8Zb98mvobovx7Mniiki4a28uL5Mxk1U9XgPYyhIy5rNkHbUqNHXeuxas
zoFMuxn9wAaiXSWYpTkJopgoUxq7rCp+Pu0T+hZ8B++oSeJA6I47ISdfgJgCBKDjWZgXcq8++Tw9
2gzAFaBb04+Gql1+xd+86+iGVI2HAVx3Dv5rDHxgAJL1if+UovZWvUW4bTwpA0yvTkFmGI7SN1mp
3Y91LoRffn5RP5fCATyfsAS8qCpkcozBYQ6iePnwquGi6vAI4lwi2WTsVjERmH8u4NCTzW9VA47N
5uzLiVSYSOFBPw+pjbhYDfoq1k7YK2+K6ovt7vSUZ5NkYPvOEmAVz2xLpLKiG5uGhMCIBOrnXgVm
SfcXxWSwtKuX4v3WGMWQvvENrKe4VNm0SZKn8SOPvn561V/vTTAfbzNQcG6Hyyz2gJJo4t7dyK2Q
4dDNght6u9yiLFljbmsvKZy704+07I9v9Wi9z/WzCtgA4wwFSxAakEN51KVrMOy8hwt/Wx//g4og
5SweffTXU7y2fKaCk8DhtW04kAlKZTjFQ2KqbPVAKlwslQmWZap/6liEdEpmuOd1iIJIfTGTxPb+
AipikNDecEXiezquBCKykXq5IKt+YjBZoBTpS9Zi11ZvQu+vkThBfiY6vh/SU96gkf2ZiNiu/a+k
ZuFChXda3/liADF5HGlyA8wxueppCVNf5bBs+oCbHPmgsdAor9zxIb90E5DPt2TfZ/ItQdxJMwHV
/qAkdZW9TH2vSdhoKpI2N/+50KCAtzYInlNftfCsi1QXY/UUwM1gCGUMOEuhnrlC8vCPspqcIS/2
Q/5S1PoCYlrwgDH+OmiBU/evedx6tQrgI8H3TKJqi508vrHQDOVrs2Ql/xXWhTatCvTjX1HlY9W8
22w5eQ1AXY2cj2GrUs7z0z2AZr/cxcGV5i9nj+0JArR+klOpq6/omgq++qajM7yTrZJvg2UbNvCm
iXGIpeMBHyOi/UmP9PejS9nWs0fqfIv0DcDn9a85wguLiz6eTA168J9PsMF3GezwNLjewHXZRO0l
BBkWB72FqLEIHo6WWW6MbNI/WY+T66WiEhZ/kdnF/54C7WZwfRnKAD+1uSL3S53eGshO2f7yeXnZ
t6R+VyH6vw3BGW3Ckncv7XN7ATgmwvHtUDkyjd2FLqjyKj4QTbau2xOVQRjHygNAff6NtnvmUcl6
Pw5JpNUDUsW83YEB5vKNdct2pgMGzWoIloHf+4lv28Nhi6k6o87bs/+oZZMgcj2AkxF5Q83WthlJ
CJk9Y7y87Te+kuDmMPEIGMF4pTy8+uJqDsk0l50o9hfudIlx62blboMO5xRMimQxg/Bw1tzuUnGF
DHfRKUyBtyt2/OcsJnJNYBS1/8AEkxkMDZ1353a/R9Z+O6H+CMZuaZAsPd0MVjTlMiIScnkNqOyp
FngrUdwSoV37k6EcDXHmJ223/9FmSqygzFBXdWgPM613qcIciMQfdlceLFjbjhM72lIZdjLg1WgR
XFCiqGLgKn4jBVAzBep/eSy6Rq5Yvu6no7PNLKYBnjRBYvrMgRWzVq0XzEPr6m7jMoYFtzwdtz0+
4Qxvp3LNo6SQ+0LUoVL1t9h52tZe30PRCTnnvzWCJi/QnqnArP/cawqKiTPV8yE/XutUd8CrvsHw
nGmulL6VWUwWKDRgqGwSUi8RUZw15lm9BQhauV4S4wJd6+MNA+T6X6HGcd8RdeqYJ01G7YywuEp7
cKNAZkgs9OxqDmQcFlGBi9o5CduE5ypokIxBixeK5pSZFXDQCM//1cRj8brsA/HOmOwidWxmwDuY
f3aZNZAwj33V3ciFQwjfgJc3ePR0SGIwjRzLAB4XeHn95uURgz7ewAPFavZD1RYWbxhiWZGoSDB8
kxHDtQgHg12XTZ7SmKe/2J6JBzIUHuW+6g6bxdhyjKbwOrKN9x7WEFusfacK3gVGjFqnzu2F3Xx1
NGaLqZl6pyi2Syl70bPZPRzsK5GPEsqALGAi5Of6dQo18shxpYSekEN5I3+Q9292tmDfJEFytHfa
2SRQXWLMJ6Xy0u0ImNEhA1RYBd6/feIAMQ9VXO3OWN7s1BC3bnFIxXcFTRX8Ek2InET7duzsrYoq
RSb1G6E1xTxdw+wCrmAkJ9aozo1u8yPiJVb2K3YE3zYvBlCo3YtNREzij6oqVoK02jEXLJ1FRc/4
cFGxWXFZEWkVp63VM08MXciPWEOha9FIvZhMiSyiyjdOM6KK6ZPJLTXwgRrDvzJlpiuNdWNnBLg9
vMBLduVDXrb4Wy2BU7Z5ReVmXM0NbeUf+MzrexzCUVW1fwJX8i2zFJ4BNXt/cvHGjevqaf0JNrvm
WL0S8YLK/h2xOZ6i0N2cO/XWYSdSuHQj5PQ5zJf0CVqQc45Ak+KZMcTtYtG9/l167Ix1Mr70bWjr
bXo5IH4s3O2laeFF/2VWeyp8VgV7PxrJdvHFF34DBejC5p2V5Gid6J89n1USw/J0Ne74bJpw1Gcz
REVwKbBsMZ0NyJTtgEnixdj1Q1Ywb/PibGoaWAsNIFdLybLaIQPenmEFAvtb5FkMFU3HBRe1IsBK
kl80uZOOpcJ+Bjsp0663tuB7fq9mvmeSQ6y23fF96K1OxMaXm23Ofd7xEyKxMeeBR0fX98SVHtG5
RR2qS0hng4z8uwhrUaDTMeRxu/P6JkxqwpGqBIDYXAtcHTfmO7Mnil5AoabFNPln01kWpjFQ6suR
Ayzo8U2QE9S6KP1fvN48/5TK5my7eq4A6qQoSQLDE93/JCwbWU0/MQDxJbqcxAkmYaRFa1J5/sd8
eIptq3SzJxt7Xb+LUVz17M+M06K8mPlNhFDYt8grihJZwcJ9HA3SfMZ//szTdmkXB1aqFs/NaYfT
Q+oOCN5KqiImU+2QsnTs6nBLA0cJlZj56xbC5eZlJrZaVDbZoPsfYZX90wbhM+jCdlGT5fMOw+ue
QbQtvVGkgcne04W8IzNslx880xxbcI2NIg2lKxJlc5xr7XAZ1DLPJucETYB5Ocs90rzLfO3eSzwd
zzMLJxIgFcsGXePzP3uDqEApup33h3gukjhHUV6jQ8p/xKi4Gz73v/BHIGQ083E5FVCJh7QF6UfI
27kxQFgOBtMRFEuYmSEQzS4AzgMwxZXYt5tfq0HPGwj+tpjgd0ZOYXgR0uLHw4OsQlJlRw5VX0by
wnq1fPC648dviz5riIiBP3qTBnmOgVZNbBtNmOPqtJdHESaVgKdgWtpogD6Fl8OdBX6QwMwhgYD5
iLx7HlNs0gw1LRaFZPs3qrcFUkeTr+5/R9Mv9p3c1cuvnwRVw+9z8mCFFSkqgdBKjU4LS94tbDLH
eUFKCcGsw9cYJrL6bOw6RdBJ7a734oVI8ytFQYDBhJRKTvmoi/sQ1UAegoxZm997wredD+fMvweK
/R4F4KBsIQkopVaXCsxwiUfj7VVmZGiLXN1MO106kVwbfBa5vOejywBbQ16777tJf/grAEIqR3e1
Fekz5AaIzzIj0x8KA+47zB3C+MrD5XDBQXhd+xR354MMZStz/1WIgqq0hzj9Pb2T9Co1G9kG06Gj
Lv83Kpo2+aZB0k21YKpoflovnrPnt5vLYbOrJ43nmjRUJ+Kv1EKy0ln0IIBWWGCTrddO7EGDGJxN
y3oqfHiFM22UNLZgnxoGfE2mVOH/QbUT8Iso04AH8Y3HGHMuoMOV82M/MX06VvTJjwzpaEinUgRe
fvZeFVxS7OKDTjQMyJKiv8GFrBtnppO8rpF+VzGPJzNl13yK/qYL8KNywqbgz4j2Ge+/L7Prqih2
6chmwo3mGm9IRSfSGPmPSJBPNaxvDIOYW9ykb3DhUYN/WZ3zWI6R+j+1VbeAn4lK7KCfosoJbX1D
RzYPv/r1bhiEt9/0YCfNXUGViNN39ykogrnbizMf9ZYBqe1L9IGI7+UTw5O8TZE9cxKux6Dry9ty
TRA/au/VVS4VV94yaiuw+GHorD4744R46gasA5FJHTtdV1QPUxoA4ICsOLzvF8WnEFuG3UCbKvDU
Zi06x7QeA8UswZGtDeIPqwbX0+BiwuHIRIMPGkbiYvosoZlsPEtOSdlyJ9Etm1eUqxCWA38bfEZF
+YTzZV9aqz8XlY2hxvOL68e+2BWtxFL+Te/IYyhCL0id9GI+2RmsFQS64M3Wfi3AXwUJuNyKlcpB
bA26fi0s2xAlaOenOqqHqnzgZTt+gBxJXFMCJDGL0RAURTveWsZkFMvjF+XxVkAkjpvN+5ryPn1P
8fApuem1csVYrB4X7oD6pl1qIU22UBYLRdo23bffpvoeTpPmimj/I0m/AdXs7yX5j+s84D7JgYzI
ZhriXsLAmPDbwConbES3glcDxUJtSozLSVb0iU2r9d/kX16DoElI8OO5ZVmsnUT1htrPxSrWjwDr
RnpGpvjT1CljFsOgzuz6GDDTA32cUA9+BV647KtpDLrKkSxxk0VNe/gUv0dqKCd7sX1DSO9PMoDI
4nKMJLVuq6z8SsgqxI0UmaadkpOa/tjSum/Gp97RGLfS2fS0l6GPR6iYWCT/GA1ai3uoDek1wvBM
zaqjXdmrlZXQbvsDvswB6XWWe4ABic9dhlV0HLv6p8JJGGIH/M/GoWOGQo/drEZl1px4ou5fYANb
Vy3qDt6Imw/I0/hwUIWPKrNJgI6H4xncKy53v/RMFdzNSZOg9IFzczC53IYIw3WKkmPJ+huFn36a
qbv8j6oTPa9qVLCmn/yj1ZaUFdRXAui9OUZhv7IxQUBeLufEI3F8iKtGypUPkFnUwJivnxEUDeBG
3zFAlDBS2+Zpoyq101RpwUir81gU5xpYmoC9Kp/mx2K7bLFQAnI90lVdpqKLDzItZOCbv/ifhzrT
eRstDtHGmFGSqL9Y9XbgexnpeTPGw88vWXTD4J1JynDzK/MT/tPF/mTKvED7u2keN7inIwtsWzBl
AlpKPqLUF1XBKgPEkmPrzSrkHoDHJfF+OjfQQM7XIn28naK2Gn7x8C8x5LjiciM5gxJLWQFUmzer
6QGm1/LQGVEDrMIotvQ3GdvuB2xMPkiuptseQxWX88G7q7cCJXKnmpSUx/GKiluAifR08dM2cQPs
lKdO7PK4X6Eds48geS8wyJxLRM+2hy6t82WnaODdOWvJcmery7dawa8oH1XzY/P8fkD1AIA4+0OQ
kM+K4Y0CykXpTAIbemTZlCLSIkzGxlcVBLzEXp5QZp9WLD6zGxAPfSra3C8Y4F1xBEcmPL6cwa1q
mhXGS6BEI3zoE9+NhPAnxLlpGWwhisOa8U2yAYWpTcer8RHOCqqbTcaWd4v2MJJV+uTeDlDADQzy
UlXMI4IeVbESiUPSDxCU2yIxRXBaLAUfem12+o3nIIBxnNU3r1ldpYKgMD7K6hptKE7qPZ8TRRZH
w0invnvgoA1LSS3IuqEWMXfQHxZeHZZqMZNoX7b19lQf9KuNhANNOLjNaxZVQNE1sTv+XFDvB25/
sHAqlCK7wXMKG6P3ZFN2vEsyZQVxrUtBFiSI0wC4A54ARndlB1y1JLR36rWJyz2AxlwSsiEWNHQo
T1DQCd5B+V9ioTHWsNzUvHEwJllbnwifR7lrHJfTWHsRMoHptz7734t8Faqs6cL6stxGoGcbC7UF
2Ofc/lIFUXgMCeCJUuJji5uyWJh/il86Cr7iOuNHzjmtV0Wi35jQh1LInXD9mZ+I8kJ4Rd5B8ssU
uXCr/j8C0lK4pIbBK5DMokrUHUSZy/c46D2HVaYY3T+WLKtt4j+xHrAutcUK1azw6B/2IzCm8DfL
HaU+99PtKyVNbjeAee2YfCfgxRtdiZL9K2OMxaE+RvBNT5KbdNIRGUvp1lz/bGldtXKE8sDt7sg7
7EkXfOLeWBOm/ZmEfFu5OdwkR0vWxcH8TVOjTIWRBscmluJVZEd2fTNij8QbgEuuyRykyYr81c09
mPANf/9+X2FJonsaFxUzPEWItSz0WqThA/GlZQk2s1/DgbzrCgD9ccqCkZADBLk5aCy0srR4htGX
yhlk55EsiiFx9x4YHWM9D+SfS65WmKHCfVV3Ri87kJtjFPkJIBFDOt5PUN20h7rwGWI0JxvvvdJY
9zk+UFTiWNcpPfbSqYJmJmJhSeDYGaznO7py9R3cg8P/LzfqL9cugpDz8qVoLZ03vK2g0M8mK+Ms
fhF5DkdEuaCOx4U7oYzh1reFf+lPoiJk5X4e+H/+3iLbFya9+szqTswP2CNcr2AhdV/5n4mTMOxk
ID9pIFKS8PUrq4FLIpb+71SWpl104gpUZj8qo7N/HdcfidsBVPCoT+uh8GuLQ/TnWoBAPqSshu76
kW24h4ME4Ew+RKUPNI1eYhUNHItnU1krKgsSkV8sEvO8FP3se6qhLGu5jxxCNEbSrMfGLX89EBOh
NyVsNXMhdNhg9hiCnKhIplVXaFviQYJ+CrKh2uMV03LQZyhQLRhqQ53xFYIg3pgjk/UHXVzUMXbN
UMiaOBTeItUR4ZJX09fneMlrXYGWCIxLz4DbxASk+jT6jMe4rVgUMgto2JZYjzD1Ye1LTVV9tkfx
RjdqPVfvqNT+It67sfbZd1qEWln0f9kMuXe6n87Dfr4vfGht+VyKXWZHcDe6j4EBPmHhQoMKokG/
fT4/1/7M4JSHX7+CfquYaOSAb7GD9slUIae3GAwSzYpgeuNrUE/uRVY+cq/iwfTnQay+hsHl+FP6
Vmfm3F6x8cuMBVYgXJlW6gNtzKuZjK7llBF/A48VmFBjkQhGWgVUmBo0MIO6YELJ0DK1o6jR0oDP
d7puEkouyS29a2Iw0YS3o3bmS2cQ+TtdfIzqElFtptAPX4lEsNiOKR+awHRpamWuEWZrGDB/eBQ9
4kqcRdvB6ltMfzaPs658ajDUO2Lyk4Gnsw2pRTmeJfGIhmu1tRjs+hPzjOjiOqBAUX0cDDNri/hC
u0bjcriphPpfM6SW6LyHLeAEx095N0avPfTIm8YqLCrwPAT+xJ3f/BmFYTOYIIZXqd9/LCAGH8n8
6Z1Git07EUFhjerJQ0iFdufTYCbLDKGdZ0a9gehNaF+iM77vgymEJzIM+jY4XJsqvbEHFbpPff9o
pfuBNohsdJ/Y6Jaj7Ex6ES5bB0Tv+wf2X0SKLQibqWaAusxsO7kuOrKUJYmQAkrJM2YP8HL5NQnx
cxh0Ijk7UonpWAf35deNfDJzFQSyCFehQhhnFOYv9AZtNajAUmpURXtuNz6KPacIko2W5QDzYVSl
YhvJjzHxJwVQ4yZzUeMjT6I5NppbAQ1Hy6U2bon66Fq7G9OzkUrdp0edIQW/Vq5/HRtzD3AqOj7y
IIsX9USHwtYx6s5vwt71N32C3Nee59fKvd/SCrRmUPoFU4Y0VZ7aIOCzB/Ex/95GqOiHJ5JWQf4H
I2OJpOnekAcxPSZzx7dskJxBEDMhCefcuwFnu6QpLXkKQDjKVIx7wnGl9Af6
`protect end_protected
