��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��,�y�}�ǰ�=4d�H���`I"��W�`r���T:tB�T4D�m�)�	1��I�t��
��8(�8t>s)ו�."[�漆���]�~�]��;�O(1#5���D���d3�q	��9/�I�w`W?ދ�S"K7��5�,l��C���
@E=D��!
����荾Z�V�h��c,Dt��&�����]4w9K_9O�=l�uE�w����[R�\�zÚ�-J�$����åCj�[�
����T=���K���h�����,������#�z~��?�G���B�~֨1)��k��yq�$/ju�YA9��SX�{@��mWt������w�F��r���������O)�mC�&�����$��^_��|�����=������A���_"�s���50��-�ݡ��kVE~�cu��'Ah%�����v2ݲK:|�g���7/��=Q�u�~��qC���
qSa�a�n�m(�]�h-�FK�]�Z<��K�b�s��'�����C$Yכֿ��h|�[@lXJ�*Qm?�аR��(�v�vlr�j)ڦ��0p�s�bv��jy�-����(��N�vהS��Y�n)!��\|9��;#�o:�#��9|TWL��L2=�'���$ƫ���19�?�:H�A���T秧���,rJ$�p}�a�ڡ�rn#9���~�1e�[e���!������{�T�7���O�z�������쉎�<o�j��D�7��lS�ƃ���F�V�:¦?�,�:4I~P�o6����2
�ԫ�#��G롔�qH���'> x������>I�nN1.�yφ�V�ǹW�)��	�3���k��c�Rw�buRA�8����\��L+p�����U�|4�}��3w���n��B�2�Y��Bر�An;|ܿM�MT�[�=��Kv^��L�`.���kS� z@���Y�'j����@ڑ�Z��1\֜;���z{�ړO_�C��m��UW�˯�1\���-�P�DE��`���_Z��6��c���꺣���ĩ��~ר�-�L6�ɜ|�S[�/h ⲳ�a�2;N��.�J	]� KG\�>oS�0_�o�C�͜�R��j�	�C�+�Z��؈���"�	���� F^�U�3���dB"���.�v�V��y8j� ��#Zݛ��ꍻ�Mb[YL 4�N��HHįt^y��Ɗ�<�ë �!�Utޕ��C��HT�^$��.�yP.��µ���$<��Os�`��A�&�F�t�P轫�������:))��oK����[_�o�U�+��{L6�z0矬�Z��y8b`��_f<[Y���ׯ�r��Z8���R�`mmǓ'_dq��G��\״���^�\�TC���~���q�����8�%����{/1����o���Q��Q���OAI�ւp�_�p�]�u�%�
]K�>�¹S��U;�(M��-7�%�Z�~�N��<f�Z����N9���Y�i`-���Y@N8"a����w�p1R&���J�,��=M~�%�$�*����e�4��^Sqx����'�@��ej��t�w(���0:��Vx�B�}�9's�iJL��b��P�����`:T	�y��W��ǰ�H+ ��z)X ��d��N�5�co����y�^Zu�_h7|F���ml��>�cb�LT{�9�s�lw��,T�)e���J���)?��5^�(��̯z>�/��ή�R��>f(Rc��;s�ov���X]crDm�� 7
O[����mjl�x��+w^<����1TC6��&?lT&��ylN�sB��<�PKD.�뒥o�D�ߥ�Ĝ�7���%$k�)�I|DMc���"=��������>�O�p�bb�R׏���(��	�h�6�	˙4�+��/��x��no�i?	�w7�Q�Ҫ���0�f7�c|��G��)��}�fq̸�5`&�7��:�)�8���Z���@8��z��F+D)����Z]T"� _s�N�14�4�}s<��(���e��
m��ʐsq6\�ݑg�F�d��-�6�[���\g��>��I���z*��e�qH�2�D�R�P�|�=�-0LG�C}G�"��ǨD��NЊ"���IoD���f�s�`%�v��[Rǟs�R(�>�V�F�/gN#A�,x���޻`I��}�:p�8��+�F�����Di�����1���A�PGZ���FS��:�{�k��7P��w�g�p0.��2��я=0���~[ЁUG���nM�5�{�b�|�u���VA�;|ٔJ�AW��5{=��������+�8�g?���P	�/y=�Ȭ���e�e��&z�)5�^gm5d�Q;e[�,�������M%�N?�n��^��l�Mܮ���>\w8��G �l����@y}�M!`3�a�?�h)��+$���e7��*wT(��o�&䗂�Qz�Y�EA;"7���?K1U)�E��Ͻ��?v�P�:���zb{T9olO�w�&\�+Ɂ|�X>��;=ZQ��k����0��i��xP��:��ȣ���QZ��q�W�%����YQ�6�~܂)�����+~.P	?j��*%h�8Q@ĉ��J�;�c`��z�����s�_�E��J-�
�6MԐ�U��QE�Ŀ�"O�M�x�v���9�ok`1~Ҏ���c��[[%��}'0V�z���_�AK���S���ѵn�<5QC��N�~t�[U6E��n�t��l���)O�,N��rY��w�<�(��X���	�QB���s�m ����n�`_W�Ri�����k@����0ݮ��*�:��2U����{3ɫm�/�v�V|{�T�no���h�#н��O�&,$��8㕽��v:g��g5e<��IG0,xY���d5ۑ�!� �VƊ����ȱeh}x]�<��d���к�Y�0���6�-;W��&�����jw�C��e�A�j�a=�,^�bg�� P��Y�I���x��A��)���C�Љg�.Sr��EǛ�>����m~i�B����5c�w�)#�!%]�o����xE7kC��*��������`_��$V����_������%O�s4�����Q�/�W��=���-���͝v�^�@X�$:�N��V+�v9�����(�_���	L�&"����0�aD2x7��mr����v'�7�S�T�d���������(L'�6�z����
*���$
E���P��@�,b���l�B�x��'q��ذxqI}&��w����>M���pJ=��(�Q���1�E/Y�Y���ĵ����r=��m�;y@�1B�XV\%܂W�X�yHw�Y
�j��gk����y�ʧj���'�w/�=2�u�}J-\n��R�d�� 	L������#��
��P����&�[t)Zw0k7�B�[�cJ�3������B#��L4vS
(��%k	�ki���'J�W���X�:&�.Ωv�&�4�*�馷�d���T��
���<LAfB�dFWJ;��
EP�^E�@NNKqC�f�>o�B����s�:4�>�K~r����:�����eZ覩�V��R����`�$`��BkoҰ��<�@w����2vAC�F���Saz{gy�d����OH}�-�cZerk��r�s\>����49��H$�v��y}���(He�17��9��`}��G&���v�]�!>Pa�[N+	U6�"�[ߐ!���3��?�a�嚟Xι5�R��G%
W	�a�g���G�3��Z����I�7yhM۳��#�6��]�s����5q�����1��nY��J�o5K[�i,Ź]�(����ߓ)c�}UcDĭ{I��|L��)������9�,��]p<�IE_۬��a?����EJ�xK-�y��d���jF1����,�����Fg��9dk����R/�P�=I
q�y8F]��u>c�$%.k�e�a)V���Kim=`pH����r�GK���H�����?bg�:f2v��Z�]����o۲#E��\�.3S�Ǉ$^YT}����dd~�#a������g���I+����&�1�kd��>ؿ��N>��z�X�f�ԅ���1ƕ..�cmF���v��m!����@i	��J�?8��!G��hx���ϬH����1�x#��4!=+��6�����T��)��痘	��p+b�~��j�R����*4��o�T����b�"A��"#������z/��UQۤ ��0��bZ��8�%�v����R⑼!�u���)f��<�Z_t�kN�t���7vx!�Cȸ�8��y98�g{3Ǳ���dp �c���NY�9#E'R׹�wi��h��3g�_&��U0(-�O�Ɵ'Z�8��s�y�N/�.�{�X�l��P��)f��)���3֨999Gd�h�NK;��`����6 `?�@k��W�L�l�'�w�8��KZ�	 P��C$���ifǩ2�����/nA��խ�����a4,e�_���%/C@�X�Ə�T0y���Vd�P�\��0v�/b[��,��FZ�O~��"Rf�����wñ�y�ɽ��&����@�V	���� C�:x5eW��א^�3$�Vy�5����mO�;�{}�����]��5�^��!1W]�����!{z��K:w$*�Z}���. �%�5<D�ADmq�"!����,�����a2�PM��8�?.=����T��ܷ\��M�1�]�b5�f��ы>�]�Y�m%��aǠ�t	d��.���š�xn^������Uv�aU�?;���,�W�Ҵ��L�8t�x����d�R%'�/m�b���lhW��㛜+B�`���⤣N�f��@�y�_�y�m"3��`���	���i�>d�������ǨB���{G5J�F>��hnu@�߿\���Z����6S9P06�Mn��(�ϱ րI���UL�teؒ���f������V_��a>�y��*x��1J�ZP��fV�
h+�B3AeY�I���	��R�/(B����9A"��K�m@�>Zj���$;��K��U:�������EO��w��NC��ʸ� :�lޒ.��aU�����
Xe��ߌ����O�V�;�8"~Nɏ*o�Q�`�AHE����ɔ��M�̩:����s��2�R&�t8P�����ϚA޲;�φ]� �n�g�$��f.ݍ��G|�zb֢�����$�^�D�����MΒKR�`��g����- ����`w�	O7X(z��w�U/!֨$2'�>u�x�n��1�LQSD|�Ǻ���}6�'̔ �����=M��p�1����Ê"2n��9m	#���f�T��rB�O)z�V� ��^�K�ԹȰ�4I+�~Ra�ڍ��F�m�l�0���>B����bU��l�X��i�f�Zm���@Z��]`x6\�x)��c�N���������6�M��+�����1l��R|t����8'�AϜ(�*8�"�������|Hf�~ߔ?�|�(U�cqf��8Rϟ{�k��%~���5KvM��Hs=��Tq�_�� �msȏ�tǛǠ�|�΋���i!�t����w���F����j�p�9쬴��jՠ+�+nX�XCG��)���-$:�9�y<�N�Sؾ���ta��\���c���g��1�P�?y|p���]Ø��XN�^ը���s����T�×�4�6��+[�5���d��+�;-��CE7Ic���ZUf����o��X���z�J����=s�n�G��ꫀ"'�s�0��`k���W"
�J�Q�ӥA��(����]WR�a'1c�A$�5�W%�� �:�)��C~�0�<�ڵtQ+W�� Ӛ���q-wE2J>gM�rP����n4��zr~6��	#o5��9��c�2@���t#%�`���e�/n[�0G�.�ٕ��5��J�\)�6|kC:Q\�y�v�����zSP���O����g�0ݬ��K��#=�Pn�'�]��Wp�� ި+���ӏL^%.�1����{f�'CL���B���i�>,��#�-Jƺ��E,S�_/ń\Q����`_����kO)�E���ܕb����S�q� 0)O����4/�<�H�S�)"���n�a;fe���۾�P�LD��C�Lr��� ��������B��ƹ����&W��)�}��jZ9#�ՓB<`8e�3q����!M��jt�����R�,�<l��F��a���j�XtB���Q�/&>���k�0* �]���?����AB��Q�@��2�P�ޖU�|,��}Gf�ȴ��$;i�j�P�����I�"&�R׉�f�h�3��=�7��v�m�R8~�U^�P7}��)<PZa�_�;���Ճ�J+��<��v���^F�TF�/�Y��:��!���m�#"���nS�_��oC����m]�=����Ak�{��Wm(������d�����E�������u�����4S�i�b�	�������>�b,*r�|�O�������2B�ƈ�[`w��;s���[�sJ�"���N��*�t׏�+m7��8��V1�!3nܥE�/���)7�EԓC�[�mOH ��q���!aV
��������i��ga|vc��-kp=1�Х����q����c��J
b�e?
Q2�����vY�=wu�OP�7�^r0������?6�d�������IK�.I��X�(PB���DC�}��Ӷ�V�1�d�\�t��Xs{�WG���So��{�3J�3eV�fC�ũ[%Z)r�4��z�o꪿�}�O])������!���Zl�6��CkV�9��[�z��c�Z�C3�>��l����x��(�Î�.5�%-���d�o��l-�c��
�{K���؈��Fm1��{�dEgcP�̃�Q\ w9,�F���P)w�Qt�_��]U���AĀ�k��{�����H����>�~�KW.ڃ��i��i��Q.ړ.�{�ix	W�vj��uA��������ac��Q���AiS�o!�Q�E`��\P{�^k���"������|�����˓�c���� X	q��-~��Z��E2vA����<B#�m,���e-J*�_�2i����+� ��'�#f�\�S��W�Is^��oņ oiS�G�� �.�,ժ��%B�Y� �$�L���d̝�*v!��#Q�Yl���m�{��1���F�9n��%@�{����H��a��q�a����D���}6�����z%�=@��p��1l��j�.����������{��ѓ�t/_�~I����D��H�]���J	 �-M�m�$J�'Ȟ��3�4��[���y�ıF�sq�F^�J^7i-�'��@p�tA���eJmiQ1�phuDk�$6 ؎i��ͳ�[YZ7�?��4�������tF�:�uo�օ
K|�X^����*�	A}�yZ���cx��$!�0�Cv����=H�x�~� f��hrN�)8һ/�*ى��CB���v⿿�O�jI������
�n�V��y���O;��|��L�	�j�@p= ��qz;��a&\�/ׁZX:�s�9|u�
��VO&��^��o�8yΛ���l��\������E�~�i��rźk�T�T�\�