��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���/�����Cc��<Nb��.�x{�>��0����=�����=8RLG�h+OLزV����ݗ�@��&�K��4cbXu�6@A��?��I�=��O�s=���
�S�i\��D���d3�q	��9/�I�w`W?ދ�S"K7��5�,l��C���
@E=D��!
����荾Z�V�h��c,Dt��&�����]4w9K_9O�=l�uE�w����[R�\�zÚ�-J�$����åCj�[�
����T=���K���h�����,������#�z~��?�G���B�~֨1)��k��yq�$/ju�YA9��SX�{@��mWt������w�F��r���������O)�mC�&�����$��^_��|�����=������A���_"�s���50��-�ݡ��kVE~�cu��'Ah%�����v2ݲK:|�g���7/��=Q�u�~��qC���
qSa�a�n�m(�]�h-�FK�]�Z<��K�b�s��'�����C$Yכֿ��h|�[@lXJ�*Qm?�аR��(�v�vlr�j)ڦ��0p�s�bv��jy�-����(��N�vהS��Y�n)!��\|9��;#�o:�#��9|TWL��L2=�'���$ƫ���19�?�:H�A���T秧���,rJ$�p}�a�ڡ�rn#9���~�1e�[e���!������{�T�7���O�z�������쉎�<o�j��D�7��lS�ƃ���F�V�:¦?�,�:4I~P�o6����2
�ԫ�#��G롔�qH���'> x������>I�nN1.�yφ�V�ǹW�)��	�3���k��c�Rw�buRA�8����\��L+p����rw3v�FF��8��Y��8p��s3jL&���9>��y�(r�I)ռ�:�J��. PWӺ���m8�����T�װ�uy����k5ؖ��$�\��Mr�pB6�(�i��pǞ~��>��Y��M������K�V�k7��YF��h��z�a�&1����;�$
.;1��r*Q�h?����M��j�L��I��:v:��2S!�N%��8	�VU7r���M�F>��+?�z��^}����eb��t��5�G^���\|����j��X�4��r�+u4��X��Ǎ�Ũ�aݳr�gˤ͍7嶙�Q�=���� ?8a���Cq�"�_����7�i����H��'i���҆�U�U;G�Xҟ�����U�y������{�p�9���sNy�D+�฿e_F����'|H��U2�F�c�#(q-�z}�8�R�b�k���?�Szm+Ō�i?\�>��Hθ���(�o
c�9}�M[qי%����oO+\�����n�R*�k_�(ۮ����
�^uǜ����s,��lQ��������*zq��˿?���߻�2�@&m=���ɮ4���^NT
@��}�2%�4�����7NI�?��r_�L�^+�]o�Q�ӗ�q��B���w��&�:P�M��ҙgV�S�`������d���3T�����suPV~IKښ�E`k�(�ݝF������T����V��bZwsP޻�8VR�+9�f��{�A}�[SD��ãy^�H��ٍ�05��HZ6Q�[����;RȈ�FX{�oZ��Cެ��<�q�f��	k���)P�M��@�H�Z��g�����Ԡ�1+5��>��9�bA���
-�V���W#��o�b�]i�ѿO2�stn���!m�V�_a�,)�O �WX�N��`	b^v-��<��'�g���2�~&�lv��|���2T���jZ�u�E�z���7a_��[�)'a���?��?L躗�&�H��V��$����m��� �o`��z;�	D�\A�@ӄXL�|�Ep���{�� ��^d��]X��ڿj�o��[�E�0�#�����<վ����N�%|�0��d_��"�����W#{�#��O90����ؽ{ :�����uT��1�>��V�N�� e)����M�к��r�U�/�f&ȏ�>z�����k���i�X���V\�F�dۤ)S������b�NH�(gQ��쀨עBC?�kG�J��Q��K<&@�{�`@�+�ts���8��(�j
q�;���f�0�9`GF��+O��l�d��.��|��؁�<�[����\�
�KO�վ�fk�H�J4��m��,|�	ه�;]�0Eez�1�r��)��'��gɩ�K+WB���i��6�����,k���5j7��zI�˶��+�3s�=�%ta��~�W^��p��U�p�,^�!W7x��6n��F����f^h?+�H�ۢ�]��b��D�솃�r`�نT<�>�f��Hʽw��oؿ��"y2���}i0{ع���F-�����>Uv=�'2	3�z�⾭3n 4l4U����'� '[<r��#M����k1���n3�����n�$&}癡ZZ�NK��uAN�drT����UIzn$��%���R0"kn�e�?KY#���d�}O�O$���� �X�#$�W��h�r�i"~[�7&�ɞ���?"]���P�`K_�F9�t���3:�_V�"
y�i�;�0�qU5�oO(��3eނ^߽ZLO=G�c|F����m����z����I�/�q�:�
ν��_|��(S9�~B��O���"sn� )��w�g'�4��NN 8 �e?к��#C9=�H����I����JmDSN�B]ۘ߈I~���Ƨ�N����6�hx@��V��HLt���D2(�����/q��q��b���.�S��ЂH�X:ov���h��7)˰��o���9ieKy�E����5�%ϒk<�y���9�u��OŮ?}����ӌ�el(#��I�j�+�~3�n��AC�j&6��U���U�p��S܋���w�&��r9�6{'H����p[.�L�q�E�t����>��Y\�0o����z\��[B�ю��K?W������,�P�#>����a���VB��4���uŹ�x5�x��V���S�#���u�02i?q�4�� l�Ilķ �-��4�[�9����@&��ؖ�ޕGªa5��@����zO��aǅ�I�m�wx*qQ��k/*�W`TK�7f�مF��%��~z�pI��/�T�^s	%l�4� ��q�zn�����e�e`7��u�{t�"�x�.x���İ*K��E�fe�,��y��|�jk�lm��sjH
��
D��"$����M�L�߫��)~��+'B�M�]���$�p��9��2�o5XX�f��"� }��@��z����>�`rj�]n��"��(�c�a���z2�z�_e�T���������s�J ,����|S۔(%��i�ά��g_���h�Fu��O�l,X��S�[t,�����+��؛���YCU�a:��뗺f$Ϯ�+!ȍ�_E7������U���))��2�?�r�z��/�<�7��>'ˍ�|ҝCX(P;�)4������YU�.u��eI��(�A��{h`o�"����x�g	������Q�1�߂��[��\��d���}�kB���7Hae���f���ӲU=�2y���6/Db�Ca`[ �t��:2�B��Db3��h���g���cs��z$�f�x��^!��b	T�D���'�]A;�Ś�<Խ��� ѐ��/�g���Y�Iz�o�>N���_��E'�)��*_Ѻ�o)��6��N�k�5j%��-�	�����^JŘ�1=��-�0;���L*�5�"�0P�4<ȇ�?v�̞�.6-T������,~�=&c�Q�g1Zދ��]��-�4�{g8�c�5=��:-7&#�䣏JsB���5�3�w�9���m��EB���s�V��&h͓D&�Ҟ�*rU�D�7������ ��Of[U
͔�eݛ��	���q�]��If�@尹����EvD`��a`�)Ӌa���c<Ȯ���K��W݆��d�3�!�daʤ��/х�ZM���-
h� b��\�w���dXS��Z�.>�#�8��6�%��}�HMKM0D:�U��ҋ{J��A��ٳ
���4�^���I缱Q�H�� #����G���O�MK�����HF�z�5�%�߶.S?�-�7"x�I���W����:'�jzO��s�������o����o1���[|���E8<����{��%��1`���nÃ\P����<�(�,�G,뮛VS���Rj����6�S�I�g�z'bQ�
��4w#x��Qۊ�=�'o׌G�����rf�}�Yz��́���~�o� ���S�7��CIMt�]���CҜ�h[V�%����Z�>��P�s�X��7.:�t��{G�/ڮ����ҽ���23_0"L��fÔ�M5ϸ�O���-�*�����#���2�*�;�k7�\)�i�*��Q�����'��pV��߅�0)�	��L�m=j�`^E����M Sm7��O b��lW@��7��(��]h�V
���gɢ4�Y����/�h~���KUuhl�zi�ltSn�sZ��8U\�I]/�9{���P�1l�.���Lqm6_t�{m9���$x�������!ZP?��{b�#�Dp#X�M(�0��_�
�B�G���)g���G��6��s��)�B/� �2�m����Xf+�]��Uo�n�8�*^�i��,�j�V������ݪI�<`����H��g��d�^�| ��Yl�H�����c-_��d�|
���V�.�כ���6�Z^�Ck*r������ڧ�h��@����Z�~5�K7䬳���V���{��yk`3�I|ɞ�D:���1ғOB�<�Y��ia1_ٺ��-�9����1甍*NqL_��ΒD۠�eT9�&�2�O�D���{Ң��
��we>���.�U�'��"��'����E���M  ���9�1�lƺk%r-r�b��V���r3��:ll��$8�����^Z�1���ЅI��.W*�?�nu	c>-�Fw�b��M���RYNL,��1�������fBC�?��rf"Nȱiߞl������ͽM�(N�z���ѭA.'ۈ����v6qn"Ɉ<�g���A�?/�[�?�Η{]�BP��,�ʷ�VG�F �{�3������;�ԞHt�j�K�4	wr��!��-� ��.����Q����d�V�Y�ڛ1���.��T�f�w� "���``� *�D���ޚPU@�W���2�U��R���j8b��Ѷ)L�7��=�Ү`�MT.,OM���X��cN�T��Fq�7}��mɗ�%���?u���+�����e�%�X�n�&oT8�OB%c{V���rjd����z��2��$;/)Fm?_߳�m��m�^�C��Ϩ�w�#"H>e��Ȕ|�s����m���7^x��']d�_�������.��^.��r�hp?2�I�x�v�S�z ]̉����n�`|J�T�]ݣo����Z0W‱~0j?u0�R+�"X^r�lS׃6�ugY#�NzJJH����NE���bn��F�oհ���J�t��L����	7M��K"�B�x��n�5i���l'Y��,u��mi@�xV�s�Z�Z�K����s�y�W�#�p�)���c�2������B>��:�ljg������Ĳ�Mp��?�L��k'>k�j�L��<�S��#����Ԝ"RUs$��O6M��i���#�����.yd��Ӌ2�#+�3����Tx��9<��2(���$^3Z�P��?��5|X<�9�ߍ#;|f�lq-of���Yσ�~t����:�m?r(�R;�_	Լ����a��U(LP�*�%g�'^G"�|�#MYA���?�i���rÇ�v1:!)sS��쿌�D<��D'ۓ��xb��?c�#��� ��c,����De����e�C��C���&<p٤P�W�]m�B_��n���_§U#>[�e��`�9����S����cF�9peά��l��o���㖇�47'�B�[�b�z����0�)�%��	Z.�����9re��.=���L���P���qqh<i���!LD�IR�;�
�.&U��t��	���U5�@O�$��u>q��#��1F�/F��p�J;/ �;����I��-I%�*_�x��D�?l�R[v�nSh�9�'��C뒀��0Ώ��H��JP��g�R��+v�]��<�0ʾgց�����5#��>� P#C?\6]�oݍ b�f��y;�?����U��h0ʲ��8�=΀�+�%����Eg���H�u)྽3Ad�F��/��9Lt��_�"3���s#p�)����8�V��,N�]D���fH�ʅ�1Nb�g�X�k}�~�e�-~ ����PV�B���Jn��ʣ�e7K'��N�ٜ���8F���G��d�tԤi@�W�c�}��i?�ov)�d�$܊�������ɽ39qfO�.ϋmA�&2=�<�c~��Y\V�!���w��a�H��AF VE��T�W�2_w[1���%C��k;�*��'j�������"�J�嘠��v�n��4~�eY���i��)7�K��!��`J%RLe�U�>xC���$�˙�6  ����R�uS�$D��<'�k��	]bS�u�`�+�
I8�x� ��R�C��g.��/\Y۽A�5�.Ϸ������{*E�n\��Y�#��7ݯ�ʍh��.O�9���D�(�m��	�eTp������������
��mc�Q�ٜ�YWY�E �`Z[if���Y�2�rڹ���p�%��A=p�h[����`ֱ}S;X��܄�]���U���%"�V'i�Zt3lW�w?Tww�o!5u�{�K�Q9��"�%iη1l����"�#Dѝt���nZ�����>�aK�Y�|qOY��Dh1�=#��&����,w[��=������K�?����o��cJ0NGF�L��2 V�9����z�C��[Ғ���M���m����xO4Z)J7���|��Db-����4���?8	>���o�ȷ�`��!�i��eT��JV�l:wwB�N��h0�
:oy��"g�	��	��4�	>�0mV�)�w1�M��
�����+f�.�|��H�:�k�7�^"֬{�Wt΃dt�gۉ�����H���P���h�Kzqcl�IAX��+�����y��o�z� �i�<X�2ۺ[˞���}���W}`�H�� L��;Xy�94˃��G�����s�(7�Ɇ�u�����kՏ�B�o���1I ��)�O%�ǣ2u��o��8��r���E����Dn� ����]�ŝZ�L����o��_`A��ʅrD�(�ID�n6�iܑӒ��3��a}�r� �y6�Ɓ6�"�a31�Ɲ�b]�k�J���ql���������lp�',CO���
_C�+*�p��T���m�zU��&�FO0�w7�����o#}�8����"��1wF��K��Ȓ�B�zF�?��a�>�5�i�pN�ZqI5���(���� ��3�]�����k���l� �d`�1�W@�g�����[��O @���_.Ѧ���w�Ȩ:�����O��ip1��"�0}�2�|�,�6<� t�C)��oZ�Vڸ��)�)���Y�!�����
�4�8c]gu�:]�E�a/��x�����:ڶ����_���{kJ:j_m�{��:�	�ʡ�æ��h�փ�V
�<E���N�9"r���=tPz�6���Ղ��E��Hd�����M,�yvt���l�_�x�)��?Rk��Gl��+E��/�(�B��N�J�M�|RfӲ>u?EN�z���;����������T������Ư=�n�=�Fug�cG���B��>X�e��Z�;�}�+F?�l�n���T��"?53)s�X�LK!ld�P�k�*"7VɊ�M0,��:���m/ a���pX���H ���犃5!-��tx+#>�� ŬFM����z�PD*$���/aP������ta]�i��4��GV����V�n}�8�������&qܻ�;LA�FIK�R|Vz��|�[�\"�f�r+�ئ���Z�Y��	q%�Oɻ@�1$b�pl'N�Be�Hi���Pl�s���w��1m��.��=�	��� �@�Ѱ��Ő���l���T�!��9�_JnF�~���yR�d� �Y��}4�h�?H�tTB	��e�߶[l)��x������Y�4��"b���=W2����
�q��%ܿ%���5��B_�W,�B�Ӌ�$)|F�M�V|Eep\z����	1�~f�\:�i8����� ���VDU�T���,"e�|����#�x��R��p�#�<�*��؋��Vh?���X�򞢂��^�K�YѭYC�v}]�����K�C��j�6�3�=H����ܠ��h��&jI���0~ŧ�ɾ���7��Zʸ0���0�$f>����Y��`mD�Ӕ����Qv,�A_��>��Ɋ���
���帋 ���hx�V~� W	��,]����ۘ�X�M❸4�;	s�)�KEc��2������ٰEІѿ)Dm�L�'�F_�]���S�ӆѳ��U��{&h�}����0��7���Qz�gC�A����_cHbW����i��.��)T�>Sy��k;]�����9�n��ՎL�S��i6�I�7F�>S����i�[�S�9�4%��QN�T�����V�/�b��"L��  �bRX_��G4w�%��r���rk�:��|.�{դ��e!րe1��#(�T.Ꮙ��#h�b_��`+_Nq���+�Frľ-���|WeݘX�M�-�;�io�ŧ?	>�]��ޤ��˴�3�x�G&hT� �_�O�8Q�#e���#p���\��u
������^گFSq[ǫU��`�6��z�Q`i��^DZ?����謸����%ݵ#�l?�L<g�jR"ʊ9e��Vڥp�jS�Y�be��i�ҵ�Ώؔ��*�O)8A銹�1�b9��Bj�k�=� �!��m�V"��5�ถa��d�Tq��=���vos?pr��XD��`���؞b{�U61*kLF�UWX{��p,T���� ڋ,����V��Z�J`�Q��y���CaŮ=9̌��A��{j�\���9��+�ϡ����r`7`����Jy׾^����  q�5M���L�P�w��Cʹ�#Ƞ2��ON>�\�m�1ΰ���	��G�?���_o3 Q����������D���	r��W��exr :�� �Q�B=i%'M���K�(������x�0Zh�Ķ������O��r�n��(]CRT/՛2�4c��.\�п�c ���;��w�/8�Z��u�:i)��9!�D�;��0%�A$	zÇ�oZ���.���Em��x�������D�u��6e�i��1I~��[�Ʊ�Ҁy��A$B�0�~�2[ ��:x��벣���u83�K zq�)tJ��vZ��g���Q���H���Dz]ȤCA!�I`[g���f����2��<\�"/�X��|��
�ݩ��{�[t\8ڑ`��߉8D���>��S��{�dA�l����7S��Q����5�j��K���}R�׋��Ĥ�q����~�&/��T��D�J��֭���h�����1S�^/�vᘓ��x�ľ�	���4&"p���
�Uo�Xz���nL�3�N4�l�2`�Zr	A�<y�ƌ�pFǋs^6���zҁf����}6A-G��6T�=|+4�I����ƐV�S�8Q�_��e��j�_B�PE{���Ʒ���S��h�XsrKĪ�S��$*b��-:&!klc�mJ��IA�C���`����i5l��}'q�4�{6e�J�ƍ��UB?w	� D��&�nC�(�Tn�,��⺵]�<�
�>�/\Nـ���Ew�JZW�ܡ�Pl"Oa��^�1X1ñT�X9���e�''�3�A4�P�kW,X��� �K^ڃ��Xd�. �+���di�h�ӟo�P_��ڤ�׋J�©RB���'���H�zĺ@���������=U>�R�0t~��=<��\��IV�-^�W�	��ٲ��s�S�ȍ�{�fF�G��3,�<b��?�}_(���%Ģ�6�^�qB8��J%Xv2��Ў���6ʴ����:z��qR�d��#b�f�Xo=�����1hE��S� �XR�RK��[�Cp
�3���c�y�8
�N�����Z��o7n��.'��n�2�Bҋ������c�i(F|cM:v ��'��w���3��)�G�$��8+0$��+�p�V���\[��Gc\��/�|JI��`�1��r��X��d�g|�l��{Q�l"�#S��p�'T0��(�WO�h<��1��^�'Q`�h/"�9��'mCD�K���k�Wa-()�w�m�Hq=u&_��Y��� 6�Dc>߼���d���"��v�_�ҧf���{ ��gD�{�V)�WuFΝ����5�Q�hanx&�h)��L=�(23K)V!�kDq0[��b结(��{Ş]ȕ0qaZǵ�Sd%�3[5Ƙ�O����O+=]l)E���Zbq6���
��/��h������u�ܳ>*�m���(���DrAìm^&�e� Z-"�i@e�xA��z/�EOβ+zZY�%Q��??�9+��[�%S����"@[dՃ��n�n�w�"9�m�6��2�r���� l`G��2�yKQ�Ńo)�������jk	�#-�/4F0�yM"H��D���qzօ����6]gC��xiN�]���2�s&N�β}1\ю��gnk��
[�l<�PM�hP�U��:�1�|��Ʒ�jGv�.+�ER��6yx�T��A��%]ʜv�	�Ӛ&��o�����i���h�<�L�I�(:��X���4Q�Ab�:>B4dr�%B�},I�t�J�M%���f����`y����&!���͙*���_����Dd��{x��ɂޱ����up�N>s8���Z����c�U;r��'�n1����z�U�.���b�ƆY���ׇ	��� .C�i�G�D�
��t!������󞡼�5������E��%~�uzK 5h����Sc\_U8��b�����^�kI�#ǝv�GdZQ6c�5��� 3 ��k�ٌ=ěe������y��<��t�"}[E*Q޳c�N7횜��l=}�J���dR��;~>��[i���f˃��IBDX
����UA�'�k�f������b�B�������Q��ld .w�U�"O7�X9Ig�.WT6�{���UD�R}��zQF��X&��؇|5!��4N�a����?���C�[w��$��R�tZ�s4`ՔSj���S��NŏV_Q\�Z'��ְ;9r7>WƗ�eA�v� !X�P@��U��-P+���ц~g��ү��s�w��g���B�ؐcJw!\ȏ�sh���w�Q�'��y��p���a$k��>���i����BAwl{gv��~����BZ�y �[��&x�/8T�k�^���v	�T���h bZ�iY���a�@�C.��Z�DZ 9�0��1��U�^pK�vTI%���v�I�ʰ���o]e��e5��A��R�e����I���䴎��T�������/\�P���\���I��f��&X� �7��JW�9@�ֱ�\�z�da\�O̼Z��|a)��H�����ED��B%n�q�5}��������h����:�o驠Ǐ�l�����A��:0\܌���X�6|�Q�o��H�B����
��ΘC�=<�)�������;�������%3!�L���S��K@Op�ܟ�~i�8���H-N��Q�C�"��8[��\I[|����p!N��>��������?�B��lR�S b�����<���\��:�Й�Q�3V�}�6k��3�5\���~��qG7����X;W��c�ue�b�� ��Nw��Rn���?�(��*�Π��
��Ԗ�$�kޠ�!��c����x���>��E5�d�5�+��w���x~�DS#H�f���ON��t6k>��ss�픻�}t�C�F�4�Ol��^?�3�������ޭ����z���o�w�Ѱ����wm���hX��P��J���ā�K�}�X���U�Q��k9|���}$}'���ak+eB���7q5Sy�B}ǀ�H_���nۧq1݊�D�k�p��!M�	�8��B�k��w���a���q�3ၳ5x���>�|Sَ?�gy"�:*����hȹf�>��G�� ����D�d��I��������|�MT�C�نf��o�F���Ν��\���$a�����wZ���Tj�QF�جF�� �me����|C�|�d�}��F��F%� W�㝀��r�������l�19R�p���Ć 
��E�s��֌�Z�J�y�b}tF,2����B�G��
��JqpO�RFS�3��Q(�w��_���-c����s�gj9�	{2��˾n�*�j��w��km;)W�=�_�Ú D��@>�� �+�2s��ޔب��/����`O' �9�x�=�G����%Ddy� W
v����D �P�Ϸ�G�9�
�9���"����W���<:{���4v�}lDr:2ٓ~+��������$N���n��»M}���9�����E��'5�.�n5xS`�k��mX���x �TU�^]@������;o�P3�F��'�_��z[���9��e����!�NW����]!���ބ�w��S幒�9@u��Xr�"t5���T�Eͣj0#K�W	��)�+rA��wn��7��p<�D��vz�&���d�	�HEeu�:�e��;��Q��5�8�g
��ܱ=.[���M�<¾J�yK�Gwq�|X�u�\Ĺ����0@7>|�2�H �ҦS�=%�QV�ҹ9�M�Ru#>q�ivSɂ�5�^�K��i����*�w�����B/��� ۑB����1�8� ��ʟ�͆LnU�,��}���&:�4Q�A ����op8�����BD�{�xR�s�S�;GP�Y�O�aK����[(�`C��(��]]	�beJ���a�t!���}�{����e9���=�{��X�}�x�Bԁ���3ElV����l��]\]�s��w�+h�i�'xJ9�Xj��V��bc�ā�9 Q��E7�����FͿ:�cJK��N�&+�W���:ž'�a|�Y�q���� ��˼P��j��P��������o:K~mQ�@�S�=�x8���t�*�"�_����-h-,�TP\�yD[�&��y��my��W��.�Ś�-���)p}��+���$�~�X���K|��p#��6#4ߋ�?ǆX�R/�G �?A�n$�[)ԭ��\�Ɛ�eh|o�V���vn�|�ٿ{	q"�wN	I\(^�i���!�g�H�}�].woH�w���itmŌ����iI����g.�LG� *��ZH3��+�[<�;.���<3��h_`f�"�va��M��o|��q�[������w8?��v�8s#=F$Ȱj��<.JS1U�0�{��e&s�ٸԷ&�9�g)��hw�����<�+l��_���Y�"<�TՂM���ʝ�%�^L ��ۘ/��Uc{�r-�'&#0�Q�P)ѝ��Mt=*+�2 f�#�%��{!�hle(�c���"���@�;�?7|%�J�`�F'�L�ݨ�ͪ��i97����dr�����M���ɺ���'p���3�Գ���V.�p�	\s��&/2��={8!���蟝]6�:,�{$'����Y�C���b2����s�{������8Y<�7�o�һ��z���`��fB�g	 s��8�Q&�����x�Ij\=N7��Tc[�8�\�H"����8g�ų��̽�o�R�Z��
	�ʃk���) �KIX�P8(#�^�v�J�3֐I���F���}�{�����b��� �7	V~���
��غ�\����Q�
O\�I�n�A�6��
Kz��=�H� =4,�QiWn\�����b@[����ۉ�D�b|艹�Tp��	r�L�#�5�\���fU!T�3�o�.�XP���+3��-۶ju�){ey���(��-Yq_�C-)*AHF�8!��p5f�*�:�X�z5��E& ��lR8���^�(�=AMK��ŷ�9�Q�ߍ�3#�T���e"喷5<�]�)��hs.��]1�m�+��Of������NxI�)�����s�"|vR�~��/�C�[D��t�C�}������dvG!El�IL��yP^ƙ]ڂ��49�ͩ��'��9�J���}1G���y�'t�gt�f��y�u-\�<�)e˼7a }��^
>L�����y����
;Q@������B%`�i��|��,kD�C�I<���9��'��%��4�P7Eѷh^��V�g0�d[w�љ��)�Q�pm�����?Op�36[H��@�_O��W���d�������|��-�+|�	<��
h��EjL��_;���Ufj���߿����/E�lcbǞ�idӋ(A��E��.SZ���Շ2jJc[�	
q��[���ƈ� t�'��C�!?�7�lx�������U���o�N��CE����m���GO�-[�^��Oрk5�{��[��XI�8|Ň�xI���@���q�?ƭh�mX��Nm5���LC{;�-<���dN�m?A��KW� V	�+�y�!h���q��4��N�:��M�k������m�����ܳ"})�'�Lr�.���H���]3p]��V(	.ۻ�]��MC'&+���R�����vw�>�u>�ZFHxQ����	�K\��=Ig�p��:s���>�0c�o��B�jsթ�W=�?�=<�<S\q������0�XN��7��}���@}U��� r��W5l�v���i���c��ydg�>E�$:�ŏ>X��[��4�iZ��y��_k�?��z�s%~*��1��^��Z�=����79Lm>]l��2x�LF�jm������Ѐ��Hy�z��G`�#UtHZ"�J�C�����K���U�e�o~c+t�a�B�����6�Һ,P�(�ThS�F6[q"rG�C����5��(���]����A�eӮ��p��Tn��څ�$�En����g�M���2��#C�e�lT��w0�Ǧ��)ępO�jU_�%�����>�