��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����N~@#�k�0!����+��=L���0�ԴZ�2�Mc���ZO�����=�����վ�	"cqw��a��TS[��{=:�����K��-�մ�(��k��N�-� 偙O��QZ��~rL'�x[�i,mׇp���O�I43��4d�,�H�����SN��d���3���r��m���̨T�I;uj2Y� Er�*p�Q$Gm���p�V�`�2^���,hz�<p��l�Bxt�5��s��\yq���#�@W���f:m��T�	,*�񞭋����_��㧋l�	�\�:��uGd��PǷ��N�I��_����Tuv� ���us�(H�~�{2H�:Zor�Q	#%�3ˠ!��iS��95�,?�.���/�F�i{#���Tp5����Ҥ0{%���2vpn���X�����@l����3dc�ק�3	�Ed&3�ZN O���z��s�yxӡt��v*}ԫy nj#��lc��m戭k[��5)�A#�����8�!�]�Z�s�M���t��w�!��'ÒE�rv��Ϝ�c@<U��\tq+��&|�&X1)C�����r�A~��B�&�����s�:n{p��͠R�X⺂L^��R����c���f��J^?��ܣR�O 1�rV���:��T�4���AD����˩�F�w��)Dm�O�b,�a���1$��c��7t[i2>�ޔ0,S���󧇳Ϟ�ᒨ�-��}�!6��Jyv�醊�^_�(�H�(y^����o#����X��3-�k\8�M�T�"`R�DF6ȕ� �,5�;Ҭ C�k���1\������k�t־9�}���� ���QHF��"��t�9 ?��{E_�7��!����](�S��0�q��w�9��=�i]�1�GʦȪc�W�XC�|�$��}q�6����zf(����լml�dz������*�eLD�*�,�m�]ہ6����D�Gw� �g��' A���FX��\өܹ&�6�h�Ð�$�(+��埧��= Eza ��찠pr[�c&��nP��x�2�TK�M�V���3Y4vIR\������ɭ�1՟?4�_y�y+����ƄJMm����@����m�����c�t�����:ud�Q�����T4���QxBŎ��\o���t�*Z�$�*7<�t~eP/`lfhg��6��[nn��#<����n�D:� ����4����.��RYF+�3��x�5���r���.��r	����h�+;֒�4d~�3�{��Ey6�r(c�d�k`ܒ1u�g��E��ծ�?��"��J�a�ċ#���VL���ҵ��ۀ�Ija�a�P���-�R�g�$�`��;v|a<��#Xa�����Vq&��C�'�P�%�e�6��)�V�0��D��zr�a���o��<:�z.\����\��ͤ���|ƚ�����_�,� �m%rW���Z�*G����Čzz��Vn;o�4�"�:�s��O��Z�I#@�u�ړ�Ac�\�Ť���F��	�L��;�����{�S�bn�=rc'`yS]�c}ɖ�$�U�P��:��s�뎲��.�e�:����|�ua?�L�;�_��� ���Nz����t3~ސ�⿄:CrT��U�����CȊ���������I������
'�_�7���&���5����&���`��<v�:��"���,n�$���]+�U^<X���g��L;� �	YC���e/GQ�^��O&�P�K�'�%(~U��
����X+�G�߲#�r �8�C� �D(�ʳx����`ܑ�y����1%���j�9�N΄�p	Js�L*�2�XB���r)�M�.����o�TZa�W�`#5�d�j��s�.*d��P�;��N}4�w��M�=pz��(�p�z�ۡ��澨���MԴ`z�}���'��r#
��Y��Ӌ	���񒽁�Ǳܮv��i��7OZ��r��F?�:F�yiFf󹺚Xp;f,�Dtr���fhe<{���	@�v��/0���O2�v�s
���*Bw���_�?X�`��[U���W:���I�9b#�VGn������f.��hF:��ܼv<��^�Y�.9E��!�Y�!$ᱶk�WrP��E�D�y<�b��Pb�}�C�+<�P����hQ#&����K��j |�=�V`�.d���O�+�g�Ց�-kg]�R����n>��?GaVM�R��ۡ�̟��b���y�4;ʚ6��I�D�J�)��#�(Y�Q����kF��_�����DN�
�a�5lou�8�q�BB�?��簖�	�E䔜���jBR-�W���1b���Ϳlud�XhĦ�+�%^�g�/��{���a�U��QLh������J�Z��6�I<$��+�B��uw�r���F���G�}k�����f�D����1�YcZx�� ����>�W9!�0�9P�sQ�����v�]uw�&2�U�yU��Xr��urRI�S��N'T:E2�Tv�;�YĒR�Y��ŝBe�I��5����2���'�>�������x{3{;B�yt�_�۔'c��jj�\h�/@a�<�>��}�w��l�ҙ�Bl�Z��;Ղ;�X��Ta�>�(�!��~Pi3`�Z�ޯy�̎x�ǵK�0p������z?�F�`Q��{&���#��VN�~�㧶X%�\ԕ�[�܆��XO��S���D��{�B�w������4��b*�b@	 �r�K+�B%�������bX�$�ҩH<���}����L�8r?�P+��Z�Kg��Y1(8a���p_�h��b(Jځ�
�q��쉉,6(uSB��c�!���`UQxC𾛧^��J�w�h;�{6<����!zX2j��Irvǈq���a]�~�.�bn�[MN� bQ��~�}���j�pA�Bwz6���ò/�S]ma��\a�S�u�=$I�F/��nlܗԃ?r�X�J-�`>���Ǳ��L�Y��1l��/�}�!���t�V��dx-e�"�"y"�( �E���rLŻ]'Cʏ�