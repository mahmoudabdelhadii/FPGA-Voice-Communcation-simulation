��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��,�y�}�ǰ�=4d�H���`I"��W�`r���T:tB�T4D�m�)�	1��I�t��
��8(�8t>s)ו�."[�漆���]�~�]��;�O(1#5�-� 偙O��QZ��~rL'�x[�i,mׇp���O�I43��4d�,�H�����SN��d���3���r��m���̨T�I;uj2Y� Er�*p�Q$Gm���p�V�`�2^���,hz�<p��l�Bxt�5��s��\yq���#�@W���f:m��T�	,*�񞭋����_��㧋l�	�\�:��uGd��PǷ��N�I��_����Tuv� ���us�(H�~�{2H�:Zor�Q	#%�3ˠ!��iS��95�,?�.���/�F�i{#���Tp5����Ҥ0{%���2vpn���X�����@l����3dc�ק�3	�Ed&3�ZN O���z��s�yxӡt��v*}ԫy nj#��lc��m戭k[��5)�A#�����8�!�]�Z�s�M���t��w�!��'ÒE�rv��Ϝ�c@<U��\tq+��&|�&X1)C�����r�A~��B�&�����s�:n{p��͠R�X⺂L^��R����c���f��J^?��ܣR�O 1�rV���:��T�4���AD����˩�F�w��)Dm�O�b,�a���1$��c��7t[i2>�ޔ0,S���󧇳Ϟ�ᒨ�-��}�!6��Jyv�醊�^_�(�H�(y^����o#����X��3-�k\8�M�T�"`R�DF6ȕ� �,5�;Ҭ C�k���1\������k�t־9�}���� ���QHF��"��t�9 ?��{E_�7��!����](�S��0�q��w�9��=�i]�1�GʦȪc�W�XC�|�$��}q�6����zf(����լml�dz������*�eLD�*�,�m�]ہ6����D�Gw� �g��' A��)�m���b��ӎ���o�6ūvO��=�W�������}��	����z
��z�&�P�K#�^Qץ�_������&�)�ٺ���/��U���WX�wK³��4�d{B9/��&�	�d �Y ����6��-�X��o0O6K�-آ6�F�,H+B�*�5	��~��6�q�?T8F��Ýt��_Kf��b�Myz}���%�l���)�|��za�ӗ*���>Tk��EU�[��2�Lu�uU��=��L��Vn����$a�9�f~U=w��h�l��r�7eg�1���$��=?	)�Q��^��(�OɦǤѲu����u�r\QD��q�/�Z�/�uZ�!���KĻX���ɫ���X�����9d_p����g\��9hӍv�d&�����p���Nh��L����+3�z�w�����N�%���v�����7XrJ6=�(���9'_��_��!(�8�}�̎~ N�J �Ky@e^^���ށ^�$�`�Ē�p���R%��h���2�ۑe��=�'�� %����P�V`đ8���]��)|\�g!��N8��-*���I����BO�<Ft��9w��(h��[��Z���t)�x��;I^��I:W���Y]6��ek�x��k�5��S
����@��Єޯ�����S|y�_�mK���k[�eMZ�Ð��0A�2I߃��b�9��ƛuE�7�]����G䎱>�P~��d�,����3�8����5���O֕l�L����eD�u�.���;{�6.)��g|�Sy�RS8V�#F���)}2KZ����� D+}��a���nz����F�� �g���B �e���:^��0^fQ a��,~�옃�����M��_�D� )��2���Q#�Oxp���w쳍�>���vf+~� ��o�k���X�5*B��J�����V��Vs��A��"���h�+7V����Q2}��81�?4�Y<�죻/l��@�~lT�τň��A'��m�8H�tE���נ;�Y�x5�Z%\z ����2��נ���X�K�����S�e!$�z1��VV7|u2>�:d��BۧLT�G�=�Uf���C�9J�w�Z?�B.$�s�K�m���"��Ɛ�ܑ���X��W@�5~�;k��n�!@]�$��kh|=��o�P�i5\�ԭm3�d����a����4�=/ڱ��'��	�L��r�JQ��ɮg=�m�:R�T���6WQ�Xæ�R���4��Ƣ}׭NR�?S�!�C��-��%�x��Nǆf��!����_q�~��xkdA���Z�W��&f���@�1�
l��O��n�ٺR>�����H[ b
Ʉ�I:QΈ"˒1%�n�1@nyHT�a����]�f`B*"�8lf�.�47�: >BG�ׇ�rݬe���~k���0���PѦ��p����@�]w��9�t�I����gEfH/�Ԡ�SC�|7�:�N�t�Ɨ_H��_�*m���1�
��3aX�R�ea�G�N!B��k#	��[Aj3�Q����Xv���@�Uޞ��'n���AY��*oB��ϓ�*��n�l �������gS�����c1�8���7~;F��IP)Y�i�/�oLG�O��^e�}��b�͏)�/�.�Zn�;W��2o�0B�y�M�ݵ�� ħX���a$.��&@ȫ��N���V$h���I�̦��I��5�j���E�U��8bq��`�
��I���/	��[)����n"CvcU!���ہ$	�ò� )�s�>_�I9	g�h���Ԉė�����j�j��Oq=��l��טݷ��S���/���j�s%'5��� �#{?{��C�c�r�Yn�>U�����������k Q�ͤ���Ɋ��,曊n���d��W�B���yŗ��D3�7�0���p���@od\|>���N��w!7���C���� �V��p/T�5��E�K�ʺ~rb.\ �]�!/��Jh�Q>I��մ��r����k��P$������� ���^�ۚ!5�P���cW{d&��aJ�[Q���t�6겯�0(��|V�&�L?K��׬�9	�>�ͮ�u�q�zZ٧(�{d2Xz
a�u�p�e����&|A%�jGi�k���S��������-�c���,�����X� m�p�r���+��z���b����8P���C*/�j����9����w#C��T�a�K>Z��j[&�a��^E�^��sF��XȀ-+D�ޝ��
�N8�8���>��M�F��=�����Z r�*� �\��A!��:�b��6�x���J0<�� �@�·Z��t�����( /�5�[6�TS�
R��>n�9p)��))wf��FδHb%�,�t����ݨ��\����|o��F�`�&������{�g�k���k����={��z�pfR��T7�S�X��}�seײ�i ���hG���T�R���P�n�2�+=�H^�>�}.��Um�/������uJv-�>���݌؃/��A<S��R�i�yXZL꽠'tB�B��&Z�����s���^;Fm�\lke_}L���Bo��a�T]�1���[=՗�n�6N��ȵǫ�l���������[��}T�8����ʓ��w�<�e,<�A;�$g�ǹ���s��3u'�ۆ&�)p�n���1�+����-o�G��ARʈ��%�8���uX�s�U;%ǌw���րo?��3�V����o��g��)Y�J��Z�}څ7�p%�όѲEk��u[=`|(��ۨ�� `{�^�|�F���J�J�pJ�(%��I�h�p�'�{����]c�������S�d�>�ٞכֿ�a�_|rB�ZR�Q�����!9P��F��"kR�(ዖ��y�-�Ȗr�_fː|/���CD�(k$�e��>��4�=ZpI�s�)�-�#��@�2�C��e�3��#�ڶ�Jt���_��l����!;6\m��F_�	��w��N��qq_8���q/֚0�{������� �ta�H��BTU�Ɯ*��W��G�+,�ubEF�z�,*��ZRV2���&p�>ƀ7�Z�g��6�ȥ}���L�@��=/�`��b^�G�}�X���DJM�M�A2[biP�Q�u�C����������@,�n�j�)�6?�>��2+��/#z�U�xo|��\���4�|�Q��QVg��E�9�y�ߺB�P���cy�F�P�.\W�,7e�\���r{H�w%_�؃j�}�d���3��(W	#��3,�F�7�t_��r�3(9�B
��ך��<}�PW�0$�0�'�T�Eφ`���3��p�Z�@V�H+����)�"um%�'�`��o���)�Y|Cs���py�^<���\��[�:x���$7c��*�/^c�ݭ"�ݟ�DTf���Ϯ�v*Ҙ�Ym��cv��e�օ��9�+�)��e[��8
�(ƧUk�. �d�Q��:Q�4c�yQ��_�4o�������1qU���;[phj�V1x����G�*��2-��p`���;<�X���I4T�{�^9��i)_��L��ĀJ�J�~gj*�`q�����~�V��q=�&U��E!�9(L\
�������+\Z_$�J9f�gW��|?�A�b!�^(��TA���N�Y�Mh��
u�!�
�v{,���������F���p2��ˍ��=(q���v�%�3]��6<�׷{=aB��������bnL�R&|��$�]��w/^LAo,�L����%5�q����a8�e)��B�U������9=�Ƀ �s;�ޣ�*�Q�W	�.���
_��@1��6�[�O��F��2���'2�glm1�?A?h����lB�ϛvM��Uø�06�%�������Śa���x?�9p���и\dG�Zm
�T���L��-!I�X�*�ؓ�}����͖`s�Z��o�9�.���M(�B���a��9S�kw
{H&�"�v;ds�=q�@>���#�������$P:�nH�u=��J�=�u�>k��0��+C�űM�}�7ƒ#�����DA)y�����z�}��.���(+:���iԿ�m���������1(���̣j;�
��&(S5�Ěq6��� �Lҥ}VneV)��ͶͰ_�1��NGG��V��#���`P[�r ��ֻ�1]
�j���	H+���=xx�;�����7�@H/,Zp7b��$؁=�
��8k~��"�˟�#���ny���ҨY�t�!_v'D�3�{��m���[�
����kѿ ��a�3E����f7�8�X���0 k�	��KU�x
��_�R����n��1���(�S�ݡ�$Kz����cRj�w?R��7�`�$f@M���μ�;�`���
%��ΐ18�d�^��e�%m��'�.�IdH
t�0� n�
�e�V2�����a��OM�e�:m��_�ޫ ����}g��n�*��B��{"��7c;��av����sF����书s�T��|���+%d���:���s�A�)�R����Ii���BR�<ǌ��h��@π������d)4Aw�U"Uְ��xR?;���b�P�����e�W� �0��w~�J����S���=̨OR׿o�����$���,�UW�1�&��R�1������Q���ۉ��� j����!^�%�
�a#[��OA	{�91���!����:�2k{��@8�1��I���,~�m �ʞޓ�Ff��;~��>e����b�E՞Co���q���]0��m<����!�ͧEVL�զ��*3�!�L��ݸEB���A��17��@��j{S�u��bi	I�_��]S֌R:M�ސ�0\�x�����b��¾�^.���CD?)� �z:��ԡڦ�2 z�����#|�u,�)0���_MD���!M�fF������]4�8[��$'�������a����h�L�l����}?ց��J�@ֻ ��Ё��5�bG�:��T�����Ϻ(R��t�D��(a��uo��[����>^wi΄;:�禥�L�>�Oʂ���P��t��VZeX��X}&.p P�.����C�������e�G5�Rg���F�^��q�����զٺ,�۵��U���
|i���x��kJn�?�I$�"����ɽ��U'���R9.ő�_����&���R��gQV*�r>�0�u~�i�EfB���q.	#�8K?�=`�L�;-������a! Rum��I����pw�܉/%�,���@��[�o�ǡ�@ܷ�/�=Co5���Р������*�'ֈ�T/m���\��
��6�!�afŨb)O�&�V��F�	3	�*��fĚ�t��%�D}&�Ʀ�ze�fc��gG|~:�:"Um���d� �`ս�kA�_[�����7�l���jE�*<W){8��z�X�Q5��J�qM#��W��!��BvJ4F��Ɏ���=(� ��Dk�YN4��v�9ї4{r�[�UP��Sל�?~�]Z �&�X�p�vU��� �?�غ��eme`���{y�֒�=,���p�x���<B�S<7G_�ur��AØ��̯ȓ��O���x R3	�E��g/�o�����Au�6�q/�	Jm��1K�|B��'�,yi�-z�.w��Z�����X���0��J?�ᓽ�qȝt���N�\�z�~y����AF6�zN������,M���~f,G��rp w��Y�P�e���nU��D�����Zs�x|������롂Y�3e��Ao�q�'����&�ԕ ���E�l(H]e�谞`w�����wQ�<�9�6��"��'3�ج�Áe�����j��.IS��RVA��qSP��ch��JNv�~'Aj�k~e�ᮡ�6��w\)F�BU�����|���9;�m$��$�����e���Z׬�L%G�7���R�����,K���ɩ���wl�h��&FfvNu��,0d۞���C�|�3�]�-�'�{V�����L(��w���B��l<��g*j
E�tR��y�A,t>�kiz��P<���ٰK�Η�s�aT@�V�YE8\�Rl]��t[���1͠�@��q���0���F�������Y6n8�����y�(T�m�T�
����y�|�
!��]�j��� �{����H��Tlm����-���蟩�-��2I����}4`+��e:�� �L�� ��Ԇ�#F�,�3��݂����O�}�-PF5�����J�4��-Ov��(:����L�(�Vt�A�����-�RW��ǉc�(JGoU*�	�FhrX#CL�YQ7I����:����(huw�鸱�_�^��s����5�|J�����i��Ҹ�O�=ȹ�_�W��D"?B��\�h� O8�E%pW����;�]�Xec��I���M�����ҷ��b���7,0�Ι�nY���&� 	�4ml.Р�s�5�Gg-��Vˠ��Tn����_蜲"���a��8�y/�4�)��x���6R3��	�Ï�ք�C��
8�mJ��j�[p��+��9^��˂ӈg&2o���/\�8d9t�<X�}�io�mnZB~]�4��= ��1۟�d��o�	�C�Z���ʝ1XD��a�F�%�N�x��CE(ge
"�CA(=�
պ^I@����1X�7'TWqK�C2g��R;���û삳2��Q%h��c�:�>1,;DPe�{�y��:=�F����2��q�ت��ƒՓ5���T��"(�싋��-9��D�c�$�o%�n�����o(Y�|���T�8Úy��ƗewZ;�SqX;Q���<�(Ҡ�F�+��!#h�i��g��+%�Zi���(�O,a�tּ�}%��|�&��tx)��Ż��<���V#v� ��J�C�%�X7��@.#v<�de�@.�� ����E���d���v`$-��P�8S�&-暴[����D�8��ܵ�)`�%t�@�G����
�\�b�<;� ��*�kQ+�u��g�N�bA�y\���|��i��ȑB##��S��y"��¦��=<�w|b�v�IŠ�~`k�˧����a9��0��IEl�%
��ӄ;�&�edm��i������]W}�K�iz}�����^b����2RՏYQ���&�^��l0G����Vc��K��xj%U��8P2�o3� �l#��>�
��M�g��9��H�$_ٹ�YV���Zm]�X�Q��)� ?p������W�=���7�C�� �%Y[�%���c��S�C[�-�}�����4]�����ڡwEZ����(�#酀�""Q�4���SO��}���<z����~���ќ���Ӫ40��5�В�Ӈ�q×m�h�B4M߬�'@�MYIy���IX��g��J�%�T�0{�I�lnhL}�$d���s�}��^�;
��0�G��GIlRAmw�Rn��Iح!�i�@���?�2Ïb����U�]˘�M�h��=��ER?��(�� 1n�c1|�a�ټu�㱡�@��K���[։#dd�E��]b�cz6ڇ���'kD����b8g,�LTX:�
K7Д���#�+�n}���I�%�ey�V�j
4�HPUqTwo@�.O��L�N�Ֆ�N3�
������)@���z{b���9	�=Z�1Ƙ�S�O��4]�0^���!2�N��êsհ�߃�け��]>��A��$*f4����壄1�L�L�#��rex�[]��N<#An�2�Y⻦����s4�2�[b�T��g�8�;�T�q(*�2ǖ��N܆.�Xkb�ӿI��ç�r��	�VZC�~��͹qV����t�+�������΃�MQIvs[��Y,G�K/v�	Z���7��̞_$�p�쬙T�Um���]���Vm6/B���Ƌ�`\�(� ��dA�U9��sdX��)?�sH�h��.�pk�@� ��GoE��f�f`RS+�g�4�հ�X�0{�8�UK�%��wZ�>�_����Rf�Gd"�!�P��?5�_�����j�O��!O�ir!>��~̨��{x k�[�`�/�[(�{;��C-�.TS���D����1��9�9����������=�<̦|K�;
I{������[,B��; iQ���rR�5��e��>�*��ֶ<��\�񞒎�5si��Di+%��?���s����t]��T�y���uו����^]W4z;���/�{7��Lg�ky�x����f��,"&m��R�Y8o�.>�߷/��AHE��u��2����G;��8�[�i$LE�!�k+G
�� �eڍ��7��_��.��B��6��p��qD��qi,ࠏ�����.1��%��ҩ���.��f�\�x1�I��1�O�T���ԅ�����?y:�`#�m=��y^'q�?-R���^���lG&$�O��,S|9���|���'��ޟ�v�Y#c�B��� ��VD^����� $ 7Ѫg�qs=�ޡ.��������+�����U��`@��u� �:h�;��us�AV�e�0֗+w�c�я�3:$isqA5�l+�tcu];o�N�Z%��oHH��^��2����A FLV�HS��Y�~h_ <u���h<��%G�4��>1��Q�߳�x1yz�|���߈xz�D�!x[# �_YX�Zs��M�I�u�p�l;����P�B�����7��?S-ek���	n'p���$pf%�M^4�z�+d��g8J�q������K���-3ǉ�$�:�3��ϖY�M$��{rd�=(6Q �@�E�}�?
����C����S�PZ(��c��s$+�d��&���jW��}C}v�g�B04~���cIżf�Q�]���[��Q��;�%D������]���[sR�����!�7V�3�כ��G��ˑU��PP��L�"ox�J��+Z}����b�1��$�R괼Eo�E�-7��6���.�F�UvM��X�V�1%`jC�D��^��kHB$�%i>���QqJ�-gb�K��A��ר(�|�|�W�����^���\F�3�k�Ջ�����1D�G�Dd^?GP��U�4V�I�m&�;P9��]���3A���+�R�Ԛx�|�`D"
��M����]l�s~=�mNx1/_Lg�=�T�#����K�8���b[t��@��7�YB�
�π�ȗ�]�k��{p+��$���/�.��!j���nuZ�[}��fHzC�!}8���A����"�럲c>v����`a�j-癎[ܺ[�uɩ7�F�*@�Hqb���$����	�_��(yy:JyL���N��^���s�ɐH��l�
?��/�MT��f_�Rm�Nَ%A])Wy6��-�!�g�&E��J��[�ozc�K@0�` O�5��L�D�ur��Ř��0X��8��,��[�B=jY��hq0@�c�8�u�ާ�҉S��z���M���`{���'�_�L-�����5zY�t�&<i#�L�:�>�.�-�髪�HeE����'*;X(�@���.E�^N'�=��8d��&���պ5mTm��D���K���{y�mGK�l��7�\4M����T�x�zM�A�v'�	�1�G�.� H8��"���5Xj�8t1�� R��u���hT���`��e��˞�D�ײ|3f�%f�e�VN®L͟#:E��@�2r����>��;y���p�[W�{����C�.�o�?��Qpw@OJ2IF��+|�<�x=�	�>��[��*_���38�<�Ƥ5�����̞嫭�@Qp�0R7�W�kh�{���ڲ�R�o��h�;�iS¦+��P#��e��?\�W�!�v�ۄ3����d�?��K`�MC�o�$��ݶ}��w���>bo�k�;�9w��d�D)��k�F�o����2�5�6���L8�� gjWѰ�<���OgnѰ�v� �-��$K�:�skK�UbMp���y��aO}��=���-���;.<��b��샚⣶?ozy��fF�BQ�	A[x��w\1V
{Kp��Ɍ�qSc砓�U҅K������h�K�&�F_X��ɐ^S��z��mnj��w�:���%�K��Ki�E�Y�<i�!m//���}���DB:#d}�Sy!����Zn�3��y�!E�J���	��v�^w�d�4��䧯[E�����s����Ĥ��6^hj�ٛ�mn��*�/Tq�E��������`W��+����V<�7;�AA��`�*a�l;,�.J����u��ww_��-��8����(-0Վ{4�C�$\�fN��o�>�����&��p��I����1j(�H�f#zѐǣ�0�����I����s���OL,N G������qD��v�|ˌ���>bN�@���j��X�S��x�G�+޷�f���*QQ3�d�0���.}No?$������U��\�@r6M�,��[`�2Hy��$a}D �˾	�v �)k`��x���fU3SA=n[l�qwf<�T�����A�k��ʓP#��zi��)	0�bLoZc@�jqu�9�B��g���AC�N��k�!�_�y
��>z��p����!��E�"n� ��n�W�'ӸŒ���P~V�CA�0��W!a���=���s-f�,ti�.0�V�=��hL�dn��	�[�Ӷ֝�t?�PN%���̙s�$SևC[�7��?��8��?	����&L���%}��{��Q���c�L��w] �o�t*��܁s�a��bo[���E��L����A |��Ri�Է�o?S5"#���{�x�/YO�,Ϛ`J��T�@�_C�D�=:ȓ̲���Zh�5	�tW��i��:!��?��7����Dql�ذ��f��4�����M4@Dw��B_����I��؜"�5��UU����~4��ə�Dh�ϱ���wwX���H��<?8v Jhc��i����Z��{���/����Y_Qog�a��z"Ra*���v?eܭ��t�&a��t8�r���1��Q~��fvЦ M��[�����ߘ_�}q�_�'xߓ���8�vե�C
ჷ��0B�I�������Q�i
��:TA�[�7`�6܄�늊�HS��r��*D��q7
�R%ЌdXpC��a��!�CٞP��U� ��-��c% ��AmWc`Pbj���	S���q�s>8$�*�J5Ԉ:M���$m�~T����jo�%n�X��@c��1!'��t[��`�W�aߋ�E�6�e��Rc$N�>I�=��Օ���1̹��ݻ�M��8P�['�V/-����I�p>=� �]�X�W"�Q�+�s.��v����b�Sn�&ͱY�u�w@M��vt�PmmA��5��1�p��s��;�F]mIo��������3dA�K�K,V��̩�;�D��y���e��CtH�ѱ�,�lb/�� E@vz�SH ��|ea�Nn�,��#aoZ^�e��X)>4]^�lӠJ�^�)�;���R�b�X&�]-��"Q�4E8���l^	0��2����R.�n�NZK��� Al���X-�ѱ�=���
�g�������WMs��^��wqk�M<c�~7�n4Y��j�,u˺z��m���	v�}^�{~J�Y��ɺ�P|a3R���#��%��_յx`a�Yv��o��<ц�%�X̧Q$❰���5dC�� �8��Ǿ��w�7W���lH��2m�ēk-���a:�J6ʯ�B��$���^���W�F�lL4qO�^���U)�oX��r�Q� U�!1�c >Qg�	��`!�K�}�����H��@E~��J���ީ �5�i^�[����&��[ +����=���3���ͧTa��@o��w�����iд�:���s�!�DB���-�oO�Oק%եet�5p� ]�S}~N�,-z�������/� Ã�ː�̸�B��|-
 C/�jj�<�5� �[�o@l$NЦa�1[
�n�<w��t(:���*F#�����W6�bP���Y�CFz΁�y��-��A�cd���t!�5�i�:=���b�ߩ  �4��\�$[P�7zg/��ނ戭�^.J�(3�b����N��$��Cԃ���X1�e�`t'wd��;�An���B��dҪ���)$&#�������-j��!��;�ޙ8��HO2!6�K%�|��PȪI��L�b/Գ������6Alr��,8k�l�wE[��?YSr���*xX`""M ������b~E(Ma<ݹa�?�v#s��B��$nBu�����鳞����&娝���t��s���d�Fw�����@���0�}�K1��(_ztA�d���A���m�yf2+����g��%��y���Ũ�ꨫӐ�V�r�0��UL�1����f�{^V*9n޼݊��H�\t:[M�����I�,�k,��#T��Ec��+��ŗ�hO���G[5�5�%�qd�z�&L�,U�Id5e�)�����'�r+���c������!=�^�'�ji� �sb�Q��(�e_�xrS�,>
6�Xw��x$)�̰�g69�߷�AԄ2�����]zHJ���\p��1�V_rT��e�y��-F�{���zp_E0);@�='�{K�;�QI�<�K�C�1����Z�m��!��i�����t��_I�"�+8œ4"[��y��B�\�7��r�2_�c�	b-S,$A�v�U��J;Y^L�Sb��>��S}� �~�1�m�H�T~�~�9�%K�rʱ�ԙ⤙F6�F�4�g����R�Q����غ�+��"n<����
�&垒���4a�O5���x�uP�F��I�Ŏ�ܻ�$;��vL.���Ŀ����u�L��)3+�H!)Q���Fׂ�
��q�yFQ��"N�Ka&m�WL|;3���0�| A��۬����\��5��ἍND�տ2��qz6鮵(��c }�Rtc�F</�>D�R+��0�@W�z(����[v�o�q8���IB��>�7����HD�= �Sɨ48�hZӦ���1k���k��U��{�ͩ"�U];��ާ�B8�E=c>M�y	I���_G�U���0�H��7�Q=g�a��N�o�IM�)&����ٷKf`�\��!^av���/��X��!x�X�=�\��V����<Y.i��5;��c�dT$�n����}k������k����r��z;iĒmU�~�86�	�L2���M�F���_�{U|]���N�b�K��»����R+o�S�e��f�,҄Aq	N|����a�=��`��j'����EX�VFkV���E-������8^�7�=�O-�b�O����<�H��-3еj��N��t�ڂPQA��H8�����������dA����3io^{No�߇d&� �,�# w�����k��Jo����I����!�Ʈ�HQ�9�5jy ��<��$�"�(r�YnBg~�p�E� c2��!�0�A����j�D��A#��hJ�k�6*�y]��u����}}.7R��Se0&.�eV��ml�r>%�
��:/Qe$L�)�	s���*Ch�F�^M�ºp�� �܆�u���o-x/p��%�OX+�G�&�Ia�c]X9��N�H-  E���9����IP15ϧ�d�����2�$+��aY�c��]��}dݦ��դ!�jHl?̥з�RJCD���^۴�5پ<<=�xٌh����<ޗ�낚ZZ�Ҝd�����;gsg��Z�k??pR�8�u����_��``)k#@��E����t����h�����V0�z�^0��u`b�|g��
iS��.�ؘ.ދ�v������x�6�B���U��'tƯ:4<��e��Iw)�pz�j��Z�����H5�;�9gc����8ᄋ����(�-�E�?�u�De��g����C;Fob�,�����Z��u�^TUcOڈ*+t�'��ZdQ�Ĝ�2VaA��`�g�i�k��y�&B��T{>��Wx�i*Lp�Q	��ףDb�������5�e�� ��d��_�?�+�q� �p<��g��2-�NA�B���C�G~)�������N��S��<,6Ưu@��Hg�IWN��F�<��y\�2��P �� �(�S��eRwe�`ǺA�.ǐ�&-�X��5�p�ی7:.	�}�n��"�F�'�࢏� C�/a�NF2��bb�@�����DY�i����}/�f�r�y�<�bӢ/s�����$��h�8cP�Mz!&�p�Ԓ�q-.pD��8f��Y<�ʪ�ob���M�8�.ћ/����i���~Ia�|ۇV��	|.�R
6�#��<���Z��V;L�h t[|�**�98F9"��k�� ���v������v���6���+�F�]Ckz�m��Oo��4DP6�\�*������ c�%4z�k��t�U��S�	��͸����I�!.P<��TB0v��<�yte����|����E���h�6�19A��Ђ��������x�����;P�(Q,~�4�g�b	����}:a�b��h	���A���'�]|�PBg�S�6%Y�2��6�қ�� �|���Ϣ��6F�q�f�l}� �j
E�&�g�aK�8�;��v�Q��˹�c�`Z�����Ɠ�B�?�u�v$��������V���x��On�#,��v�Y�����U;�?N�%�?��������'I�&��$�4^��}O��~�їz�_�\�+kX�P/��j�'�L[*HPB-}���`���5�z.����X`��$�P�%�����o�
�'�u�(�9<d��T����Қ�Ӊ����|��:X�)�ݲ�o��1���ɛE����ʖ���Z�v�s�s�A+(���TJ?;��B�����7�������9�a��K��u�"�+A�7�Oj]��yԖh;8!�ɭw�$�X+�X�R�e�+�FOS�U!���1�5�Ơ[s����ׂ%�=���y��=z��	�'L�	�?w�L�	��ײ١qY�����v�(q�?�������ҧS.��I�TyĲcà8���$@3���v��H��
4m>n�ͱ�F�9uH��V�SO�x�?ʞn<nɇ�+0V."$�?���j�t�[$����`<�W?�����wJ��[n^�׿���Ä�/B�[��q�P��
$9P,���(7E�Aŧ㚻�X���~�{7�З��m��:I	�V��h}$y*�$ t�.9�]���#��KS�7EN��B���4�(�Q�d������y�w�7Є�gxYjhz��M@1���}bI=����"���n�-TY��;r��Q18�\�`O'����d_��@�ە'܌�ȡ�i*9���E8��g�����I����w8k�1r�V���7����YEs$�d�G˷`Y���,���qt��e��2���?��ĨV��߆8h�x[��e�f��������{�9D�`���ĕ���gh?�Pu\б$��|�{$&x@qΈkq����Z�v��]��,��y��P�Ζ��@I���t*��������w��ͨdW�C��RbI`�D�X�����7��O~π`�xe���#j��Ͳ��