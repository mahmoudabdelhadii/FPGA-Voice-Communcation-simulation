��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��,�y�}�ǰ�=4d�H���`I"��W�`r���T:tB�T4D�m�)�	1��I�t��
��8(�8t>s)ו�."[�漆���]�~�]��;�O(1#5�-� 偙O��QZ��~rL'�x[�i,mׇp���O�I43��4d�,�H�����SN��d���3���r��m���̨T�I;uj2Y� Er�*p�Q$Gm���p�V�`�2^���,hz�<p��l�Bxt�5��s��\yq���#�@W���f:m��T�	,*�񞭋����_��㧋l�	�\�:��uGd��PǷ��N�I��_����Tuv� ���us�(H�~�{2H�:Zor�Q	#%�3ˠ!��iS��95�,?�.���/�F�i{#���Tp5����Ҥ0{%���2vpn���X�����@l����3dc�ק�3	�Ed&3�ZN O���z��s�yxӡt��v*}ԫy nj#��lc��m戭k[��5)�A#�����8�!�]�Z�s�M���t��w�!��'ÒE�rv��Ϝ�c@<U��\tq+��&|�&X1)C�����r�A~��B�&�����s�:n{p��͠R�X⺂L^��R����c���f��J^?��ܣR�O 1�rV���:��T�4���AD����˩�F�w��)Dm�O�b,�a���1$��c��7t[i2>�ޔ0,S���󧇳Ϟ�ᒨ�-��}�!6��Jyv�醊�^_�(�H�(y^����o#����X��3-�k\8�M�T�"`R�DF6ȕ� �,5�;Ҭ C�k���1\������k�t־9�}���� ���QHF��"��t�9 ?��{E_�7��!����](�S��0�q��w�9��=�i]�1�GʦȪc�W�XC�|�$��}q�6����zf(����լml�dz������*�eLD�*�,�m�]ہ6����D�Gw� �g��' A��)�m���b��ӎ���o�6ūvO��=�W�������}��	����z
��z�&�P�K#�^Qץ�_������&�)�ٺ�u#uD�	' �/|�qf�M&P)�tL�x�?�u�����ҽ�����*c"q/�\��YDl2n֢�vtX��Q������ǰ�6K�gVL��ο��Q�������-�˚e��"gb�_� L01�D��ثU�8-��Nw�@�$[�>V,���6�����=����{>G6��v�����φ+Y��	�d�A��b<�)��Gp���k�(�vWu����!5fQ�s�}ɘ�V�k�(�\g-*����4:`�ky����sFY0v\~��$�"t��d�n�˞��5e�*�1/�v�X��^�$/$��d�����*����=Ґ׶îƹ}��k�w�x�)L��M0j��f�E�6C/ 
v�����^��<�(��kl����ϓ��I�1~"�ւU��?Q�PG��9b�o#���W�����2�Ec�����~P3B��!+��8��b�}i�NK{����1��r{��h%� cBӈ䒦�w{�s��u�˺���I�<Uh����)c&��4�͂a)t�}\(��#$�1ڿ�r�s�F��������ikV�����R���簾��|���iO�ed�P�Q��ˑ�񬬒���d������ϢdZ�1��BV��	��7ury��/�I�Q�Y��{�㥪b0p���>�m��Hu���}�u�~[���4�W�0�$�t��--I#^X���glW�Į��i�{�m(�rZ~f �Uvj�?r���JC��8�o���]v܁��G���8<��
�0�X���\;�'	�9:V�<*�8�s�����n��G `���T�r�p���^����.�6S�I�c�	-��-� �%l`R'h�2�tmh~|��_� �to� l]�X��x-Q�+�_h#��KpWYN���Ζ��Xo�&⒕�_Pl������$��҄v6�z�bH�����#!�R*���]z���N��μ�Ls�)
���� z0�j���Bfs%�׽Dh:�Z�e�n?��:tCd�ƅM����Ҫ�.>���'����Sy�#�K&�a�f�o�l�U�Il��IS)6���餑u��{�T���f�}�z��3W_���e_ɶ�ßr
%��~��'�?jҵT�=aʺ-�"]��۶y�
����w]3",�eH����z��F�ἎQ.��3?+N�<+)��I����@(�`��KqDs?k�]��*H:��uH�豚�b"��7����a�F�i�6t�&&C���4����N�56	���X���N{TVRL�P��<��:r醚�q@If'/�Lm6օvI ��(m֝���R/�_�i`�O��{$b�>:F�iz�%)���/�i,�{ڨ��a�>܄1����+Ny�����ݡ'E
\�QbcA��'=[�����Q4{��8�=����[T\n��?=I�(X� c�a>(%������lQE�(������U!�u(�#qz!O�ہ.����6sm�?2AvPT��c��=i�$U:[L3�`����=H�']��,����zE<V��M�uD����0 ��1�����g�E���R\E$'�%K$���5Qp6��A�e��5i;�0� \�����Ǐ ��[�JaVaqlAi"P��_2�4�?! ��	x �_�f���=2�;+/�}:=dC�d��s�M0i��Lqy��A������)-��+AA:;B�c(O}�c`�+�6'*8)i|�r�M�����{�U�k��йd�;1���h�����l�|�|���;OH]� ���Fx��lҒe�M0Sص�-#Zf�I6�NR������czʽ�	�A����7��5M>�u"��Ǭ������e�TG3�� ���9fM%��b���vY����mL�%��G�@��/En�n�c}�С��q�#Y�	�?>e�h�x�{�zש�S-'�/��u�-ܕ��;B��0���C���tS,���M��m�������;j:]��-�oP��M�.��/�>��6����CA�	�"r�`6�����>t��{2�2�����>�A�@�{кD�	�1t���V��I�)����O�j��ߺ��h�����:2C��zVa��w�L�z����m�O(�,i2O�Z����1�JI�>^����IJ�h�ŗ�+�C��9
�g���U;��3����E��e��+���KШ�|��!�DVG(+4NB8�"���,tC�8�NE�A[`�b|{ٽwŜ2ykc�$oY�f�KGH'JW��Y�,q�k>R�^��A� ��~h���V�Ԓ[�	���;T��$r{�Y����/@s��/����k������~���1ĬE�y4������s���猱���]���I$���Q_�q�侟�6`@_�,����B�Z�'$�#K*3�g`e�^�+3[nK��U���5%�#G�Gt'���hm�iH"��p��"�L?�n�j%�$5i�E�;og��ͯ()fl&�����Y�7�x?�'�/�������<���˰�[��6ݡ�����|�db���p����kiN=g��"���uE���8Z���Z'�J�L���z93�h<9�� ��K�`�x���Gr�N�%�2�����	3Y�X�b�k��\n��.�>Dp|3�g2M �n9v�,��lى�-qʠK,���b��P����	�bªJ\�:�>���`�>���%ڦ8cJA��ˌ{���6Pϝ��=�����F����Ne��������5
#&�xJ���&����/Cګt���c�K�ϛ����pv�_��K�����y�q��u��*ǣ�xb��������t��1U�!�l�D��φ����^D-��)1�ބ���b���yH���MA�2����S��2�6��yBW���e� ��%2!k�������T�d�Yt�N���b��> �9eUڦ�ĭ!r�S�$$�N8�,>�����Zzȇ����$t!����j�( x�!�(�g�i蘩��m�M��I�&�0/Y���:�X�ڥE�A�qRr�d:�b���n���U,u�rVEp0�鴶=*	��o�{����j��8	4U�$j����ʈ%�!�n�U<2Q!�g�e������~�q����qr	��U={�8mh���#<�Z�mR}ʡkx��fw���@�=D�=�zqh���&�ą��F*9M���{%͞���t!fF��!̬^�~���θP�ī��h�^'TNsV>q��H�w�fck/់�]�:��p������d�ݬ�5����o���RxH*�\���n#:OrOk�B]�w�]D�
�|�{$�,kE��DZ:�yw����;aS�{�n�P�**�J���?��b�/~�-�>0^���(x8RM��rBXߢN�r���� �E-d4�ž0#u�~w0g� t�������}/�]��9��w�;]`���b�a�\�3N��ǃm�裂��<d��*����3��R���4�3u�SYf	���aL3�0��tj��z�'����w��Q����@Y���[����ק&�Al�����T�*/\]��9&*̒u �A�E�����l �Zl�����L �x�b����)��X���;�!A��������V��^�ź/��H����	����Y�{�\�*"^�h���lE����@��7I�����X˙�b���a��%_D�T̺^E=��G+�PY��a�`No��+�Pe�ӡA�2�g$K(9���e�[�SV��Ɗ
/�z5��Ӊ�syc���au}[B�pj����(��o��]"����: �m_%� ��mf+ >��L�2�^�yC�jѥ�ڑQ C���5Du�����哔]����Y�HpPC>�� ��V^�y��a�눛IK�	���+�dTϓB�W�CG1�
�����\�� 􋓽k%ZED�Y�o�M�\{yV���{�F�u�O���'��ר��\Zx�;ɷ&�?��2.��Sl��������)o��)��_��^�؏��A��Dna[�´��7��lSV�>B�h��I*CWp���W�����d��o�Af�v��lj9,���	��P}1��o��0G�;y ��Z&�b���p�qw@M@����zB��Qp�5	�m%�L���X3o�܆�	t,�6A�DÎ��=�3�^�/��cL\���J�IZ]^ڄ$TE��ɑ�#��}�0f��j۬i��2T�h���8+�g#F�����F�W������������뿎jH���t3w�pqN�ʬW6@�����h[�韋(%l����j<�	7��̕��L�=][.��r�C)T�F����X�>ڊ�1��><�&����&� �a�o IVX����I�1�o�����_[�4�ID4�&G�.��2����]�T �:#W����)ӡ���u�Jq$?�q�8���ۗ�����=����$��n�{��|�F��N[@LC-E��&���^�lN~��l<U#1�����Z��"��Q`32<bWO�J��m�o���O�{LȮ�O5�`�=�Y����(���j��[q^u�c5�=Ι���I��SQ����E��W+�!�_�9"ǆd�Φ�Ȩ�¤D�Cn�ͽ��i�!|��X��:]���hk�K���j?,J��a�zx�h�0��H
Nz8��Y.k�K)4�>���e��`o�5� dz�R:V�C|>���t�dh��2�����y��Ce����F�bJ�% X3a'�-�{�n� �r�*�	/�Rs��̆@O,K�:�#�X�R��J��_��*n�4�\��èj.ȵm˦�R7����TJ,��*|�>� ,e���� F!�]�Bt�q�T U��/;vz�_��v�sൣ�U�e�?���^�~QzC�ĹHy����5�2-uns�r��c1y��]���@yk�/z�m@1A�~R*��R�N��|��3�zQ\EEbsV�|��^_����'�l�{�=����/�,K #�!ADm���Ď�%���eׇSZ;ګLf�!碷ρ��´C2���{��'����˰߽�}�q�Q�~����?&����1�'�ϕ3��N��$aS��Q���g��