-- (C) 2001-2016 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
T1Gx4MZ2pulq3QTce+2shw49OPU20KZxZue5UITxo5q7xUFzVc9KzJzmiDU6gGDCf1IPrcRj6544
RBY7kkgGVwJ9GZKq7Sri1/E6K/xeEObsO4Urvy4RstwEX86pircbepPhoYGtT+BaEjBwjm+NY75s
Uad9jPMkQJN8m1FheovShvDnxIXSU8RB1ILcuxt+meAv3X8dA/zvwBg9tq3NI+PpytdKySNgwnHX
dpk6irWh+7L1Evj3BwHiExwP+jZhDpo5tl3PGYBw48RnDuy9hMqV9Yrmb8fxQILEky553jwJ5b88
Dr9by+mFtiivaIfGQ+Ny5Q61ug8DhBNmicUnJA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 23248)
`protect data_block
3IMmLGjSuy2fJMg+B59ihBv/8kef8XDe45xJVIR48+lLJi7lOfrzYr/Q+R3+d9RxWQBnnkxPu8tl
AyNzjtBFOO2RQLa3djxkvwXlPqeQPr8XoroeVB4kpeCSsRIEKe4pp0StCMqDpcxM5Qtn+xVqAPKS
slabvuXbTikpvNerhmIVpJYnNKNvqsL6QxKpOmNMxVh+RuZQPXRmlnWA/OvXWI15rhAKyO8Cq9i8
EOYoUa6To98B62YaqSjkBQcelxOwzoIh6w0bwrP6n1C9H8/LeLWHbQeFnU0N+EEU1tJoEVAwW14d
hGexa7oeRFQApBrTBN61RN/rVhKCeiFHYPTPzqEzybPIosjpa4xCA+NDKXM/ey+cUOL97Q+8sjFG
hwi5Hbl+VS/4tm7EPJZ7NJ0bj1s1eMIXG0hpU7OLjotDOU1vo8IdiXJv5YubabPFz0zxQsauZmIP
LT4XA+UocNnkmItEuabWVdmvKbq1WtXkx/FLOkl03mipwRSqEBLV5DfqffoTxEtQ4pY4PXIq2ReT
NxFlcOj/dmYeijIeFPE9Mqc0g+Vu4YGrGkCsTOV8Br7DvXSIoYxxJgBr+m95sVHF+5La1MoXr8Oi
vGmdBWYMO5Ntm2nka38AU+u9RpLXZDC7EBMkQze1saV6G5i+820tWczLcVp9SWC7Eh8F+ZOFrLDf
NnhHBBIPZDWK6NNlrh7RekLlcpcmPMJHmMBkI1yLKJZmmgDhig7T43PRMXUmnVnRVnsfquuVhihW
ETct7EPrD6BHYA0mz8wDsH/4SCo44BoNOkqAGDyKbXjQ+nR2ymk9YmVdPfN27l9awH9pAh4sKnoO
uEdThF1KsIx7I0IF/z3EIb/btpx8C4uBOkDGomm/hgVYX+aydngV57BQjhaVjjppHlSJvpnSqw7D
C4Ypgq9kZs3oRjL0gRzIs14dRPSZN5Rd3BaZTcFerP4axbke8D+DJbl0IZfAr+vBrwyDxLBgqD4L
ICZ5LsXZ1rWh5OmB73DDQjh+ATcVI/efYgBZuwG1uCILq6JnQ00W7SHq5iSBI9kUkCHPBtpFQXIv
HjDoNSNCwtVbZlivBLvkZLdkiXzJjE7ECKwChXRuKnOVooy+1SIi8r2/EQ5jclu/poDdpNjybIKA
uODr80t9M30JXL+vLp/kCNz0QPVt6YuAzNdiqMG4ckC5CRNvf/n9g5LZZMBe9UFVz4nQglunCKCo
K67jYVxVgCSqpMEJ2G0xn7i5clgaRYcyx0azz06/GRs6a9XPJPXWwrdoCufVL5YXtGHbBBS5nAwm
p8r8eqNuNTRa35y3Oy1m/y9aGakxLn4/4hcXaKkm5q2qTKHzus4WhzSQ5T8kpOMD7LiYgM4FwTR+
NDPIRxrHEh1nP1GAAnvOS28gPl1y9wjU1J2NiuvZcKBh3TPMNjLa/Vs8gAikHD2g+HYv1zokZTjy
Wg/MqyumvbpEJpwdU3uA/m5ATGA6B3eRdGMof48Bv+buj4XURXm9Kx1fmfAKoskhENnQGrH0eLd1
Gw+57GxLY99n2unqKzOcpa90ar2tWMPErMZzTsuFFjzSFFavxxXOLF0Q8Ah7DnLrW71618kf9zen
n4yjdg8RoZeHdl/6SrOgHzjQhIo5RxKS0Yywxgs6bEWFw1vjyDEs2PuT1s3RgDuHDM0y5tAH3E2D
4E+/RTi6sKmISghm4ze+BvBYkF5IyZ1McqTQY5VhR/c0J1VdRCm+SUsyyVm5scDx6Fq7vCEFgU3K
mbBVz8GPDbyGQpJf5HchHIZNW601wOZROD9Ddj9wEoObtbM33gUHIQQHiKBO762bhWlg0AcGrG3A
qDLEtEzwLvNGQYACDAqCQJ1I2eAnSVe0R1bD4ZvuSG0Yf8WewLb1YLowD/iZZ8aCgeLirpeL9kOw
uGE60J4pXczEM86W1nmJASXXNPjfAGiLoU7ENbxsNHvD7k0d9OxBvY2yJ/Ji1Z5JE9eUx56m6S/c
drg+M2nYH9muKdx3THr79gQxf+SivsEfChCJKac4NK5J9L1CV986OhE1yYM7enAmKPO6Sgq1TIK4
JPy8MjmiNrZ12DI+BMCW7HuGM66ppgxndwmJrTBtHKC7Lsoub77QvL2LnV8KGQz2J0cCbbNqtZT+
mzvcLSH/oJSqf6rr2n81vw5dWJ/dmix+Nl6CyfhN7w4CS/5stlsVT33iuewqaO11y74aAQxGqg1a
jmUUa1KOm5G2I/KZ7r6Umib08FDTAYOOQw0DfhcLRfrUxMp005iibBgxk6vMSm/3njvA0+aRyLRI
Qn1XCpqlKeGa8sLJY4sceLUzCKi3PcbxAvi7KMTd4sxWEKPxG38FWc2ohb6xNTJRQtY7FpD/dLft
3uufcn5blzCoLUgVR5DZNJyaYxO7nzAUmukn4I9NranWqH+9HcAwAspskYWby4klTgZl8uVlZuMX
qvVOAg//m6LQqlWIW6tzkg4hZ2l+KdjEN9f2L2BAo9c/bs+6eHdItjF4NW9Y//tt7BTq6t5y8i/F
vitvsyZ/cN9v2wt1ITFjtuZP8QA6PBgKrL2Q0XgQzWgSzX5O0o1TV6mFYwxeNA63m1QA9GwiVUg8
/ohoLQ16k/w8T87HN5jvdcjN2s7MtWf1jGVF0fto0zL9ImSuUBmm5aJysYBxag3osDh91SwGeLql
L+xRklrguK8JBlAy5d3B0IkmC5A5jId2s3mSuA0tSIQcbhP7jcZRucIegO73GoWKDH+JDeR/Eky+
iGHv398xx6TflJztVcNtWxp4QuLlp98a8gvHYZrzXIqs85yInSpkmTJMgnxcrh/jcNAsuwPK4CR2
N1iG2EyneQd3FLAbK3XnImYxTctrP3jwtIEiRtbI0fTU9ztUfUkzg+WM9tfbSVlb8XV9nBqLRluq
mEONWMdlDFMoYz+om6HePGUljEn89DcPm40uZAMBvVLhC0pVfJqzuDAslH7jpjcnqxBMVMeyrU5o
IByBoORaDSrSiHV41LNBLx8IYsTGMatfMGasrtZEd3gtTQEMFhE6aYyZEm9MrtesK/OxEAnBacIr
/cPOknA1CdbWk4QUl/QqZZZi6vFydoYvFST+1BAvTgC3WaU5WRH2h1DpQOiHmIzQTZA6ChYjtIsp
5EdhHqWRLO0aNDlxxJgMwLllo3cs373dI2WcPbaQQf7AUYtH9DPrhzUTbw5IfA7p7YEqeZrieRDA
ABDpJ7hDeo9hrsKjAC33MHX6FniZMTCl0nXiCae4r+Aii1byk1A6zvIQlOyHMllYU+t/q9dgM0Ep
jfOgY7X0f6b9dil2ToL72fkExQDrGdHk6NpQMl4gvd3M9nknYwOrp1sn4tzBDsyVLF9YFJswFhLf
Qc7nnhSFD+x+vUH1yBSLVPnFldk075pRODVX1SUPvxSz9pVhHeE3lmIL72H72tzz8cIBaNYiU5+I
9K0qMUL7MXhrWrIQrrZciS+yf8zjJly3iA4Ovg/MDxYDVoaMjbnSfGlBqEb7uFPPQCixdjoKI3Qe
MYPTWZKhz7753itGScmT1NLIoRZDPtJNUEj41Pi3tD6iUCaKbFe2iDVgCqy0MNqca6H2BnTjMk1V
iguAcYWCMYe2++HIGjaEspB03PPhSWAxCbJM1PmESTovXu530A9r/Ce0sfJXXz6+FCoABymy3VFL
+/iJkS5LA5YAK8usMuNVXz1PDmYH0ZyJDcaAOcZi52Bxw2KgI0KdoVGZsScPbhVAO3QnmmKnhVBt
Aft+dm71Y3jnfqr5MVTVhC6yN9o11fNuIgQ0oseHGYyCQlt6TqVa+OPib5KZrIXw+1fS+eVhBjnT
2vUeoESQRxiMqVC6oBLdnM0K7cBAgMt1UerpOGN9tstPIQ/fxBxgJ+HTmrsTrniSGAhXIv86oXJx
Ai29R72e5W0Q24Sswk59yHXak3S1N3BUem6TXun1oGwwbwMt50gtsTmgAqw/vBeyH4HzEjgginTo
Qg1SPlfRIiab1Abrgnt8VQIaToeePvOexraq1gUeBW5tbLyRBl/7H6j/aVT++rJQjQuZ9U+ZbBX6
TC2a/WDlNo/rn32CFs8LWuwGcgJw19QArW4jsCxowuE5V+Z4FMxU2mHKr+Ojqr0urJLW4HZXTNQL
cwfUnjv8yXV3IkOWMSJSZbLvTC2Cn52bRhMiZXDllNC+BxuxsstotOulAz9oBdoUnKTjPNKtQ42r
kHJgzA7tzmHXVTYMhF1W09K+Qv+J3CFu0c5t6GzwZFUY1fu3hHneJKW0L8qs4RvTzIVA+qg7wZgE
UaIhNyiqVltaFknMdeg/iA9dpSigJKluzIPt5d2Z+YWKGd8p5oX5x1zHEjhgvg0NvNIcPntXJ9Un
c0SLF4R5phaB2vxmvS1uyTC9OzXJZgAP23jlNvML24qFvw4QbyyTKRf64htgmPZKGuP/gEcRCEyN
+92UxNfkrg+hNiyFQz/DpAMp9cWzYAov4F3pKczEYWR1gCZ1QcMOXLftjhvUz8nchELPXpy53tEA
vkmZXiDVAlZ8i33SAbtV6Av8PlmmkW7oZWpQnXDx6GmNZaCzIYii+59bQgLHmXMyBvkFPeSdyAZG
foDtgr3iiPBF1pDakGMrUR7/VUQ6i5GOlb8RPXVtirn14k8hH2UzA+Ljj5GlkVplKG1Ow+kPMvtm
efzG6nDY4/zEGSO+ykv0SUMrDDS2/AKeTcoAayS7ubWToRAl4m+1u9KE4h8buHqiSGLO9qa+FDlM
+uPyNzzxylyF69RdGynhgGAhjTqt3TUr5pwf7DwmNxAB4LhYHI0owQt0shqVCb3AmywrUZZVZNnn
dOI4MJML2hyMayXvdZCyCE/TpIrEfeYqpIHU16dkCljcdJoH/vKDvWsbgQPsTAzAD3zYj8IAOxma
7cm946IjmcBY+5Qkv7/haRGTT236kKXR2I2xK20wg2L12tyJh9BriA7GvC/uVF2Gpc0blGt725Gf
oB/p9GNRBV3Lb9/lL9A3/ljHnVZLiBdScloItJjelAcr53W/XC3kIt6jxX4mO4S7gVRndwoLjqzX
VYT/cvUejfjgZbZ6tKhPVa08eiA0S4Mjt+o6yd7CjHiu9vqjRqG6jLTYIBCCBpZeK6IvMYj3BsWy
Rz3U9Pll86s/x2B/o6JrN2iORxJNmA+M5Qclwja/I5zXANWwO2yEJuHCyAfXWduDXnQ54i57M28M
WoSrW+ooH5zzqu6YnRI21mOUEDoynLT2OjVtGOWBu7g7H/POpwbA7aEehGce28JysHGKL31TlbiV
dXkqeHzcsFalNI/8LgRYjxB5rhvgnFfi4Q+eP7qaWvjvv0o5FB4mRIJlzB7wG9AeSu6f/8WTMUdC
RRAO1WL1zBo9mcI7XDo2iD89ZmjyMc+okHsRRsC7X2Z1/kg++imeqb2r6rppngzyA6MH/C6WkKg/
rYtXB3YWmomovG0iGB/SuQUsL3N84MDsDDhuII5xMm855ZjrtXKO8qDZFbWNKuNsSpRLexbgHxas
KfaIeG8tNelG2weUdVLuygpjPxh3sogx4Nu28aD8tH53rs0ypQ/vvEV3AeGu1BIU2A36uK/FTW0D
JbIkMfP3ms+7J2zR4R9y8SIuTgfnu3W2Urk4hfkpLfRGwuExgW4rzf8sfByfcOdYQ/a1ds0HnjEZ
YX67Ve2CY3HamyEfanLG7dhCAazB5cv+JZMu+WDH5WFaQk9dFLT27C8HZqGYE1x4ZfSP8BZE6w60
hNPfG4oSMcno8l8sSmJFkW5whU/QisaNivYHnt78TvKef059bWFH5Lsmjh1NiDb22pq35VGf2DqC
L4vQ1HJAPwJVOd8XcW6NrJ86rEPkknLXEDyC3erZYO1d1d1REa9UwtjHVFmt18eVrNJ7i85iCAFa
1rxptPu+CO43xWOQZov++zTtyGTWYQyVhOwcVafLRpWX8TOG/IE6bI5fTCa1SWv66bfj9ADcARb8
VVTV4WUNtKS+W0N3C4ezFVwDz/cu9KvsjVjKnZwT7g8DufN/FQs9EKQRrno0h4q4gedMEfCfnvS5
fFp3zZ9Ya3q+kR8Sx78ceE7HM/ncryK5c9STaQdsTqiFfOirwsEJ6D+cdazwWN2tiJR42yvcR7/F
vxO330LjFNvyIDEd8bsA3vUUskFmM3FVdLpCK3M0ps8ylCD0wM7yDBw+lUduAUq2K7KDOG0zb1eZ
LjkshcrFs/40079+e3XwliO5kKoFmOXrxxsqro0EoLRRQtBKOAr7siCGokML97h+0Q9SbQo7zVMc
RHk2FvKGYNoClNH8WmG8kDKYgxhy4zgC7MdndF28m2CdHzUSBSIu7i3m7/BWcuLVB3Dq+nmchfNv
DkWoBK/TNCfgUZ6yL0vFr2kvJK1EIgDjqocyXEV5Uwv6wNG+Ek4Ef4NL/MU/cGP5y87fLzdTCqri
DjQmgx3KA8tBXmbPpygVr+mDqRkOQfrNfEosoQbi4+4E0giqD0aswPMLkclti8BDcbMrNHi8uJsm
5M+I6I3SzMq/Ff9/6kG1b2RrtbuHJVPz1FT6QqYQvNrnQu3AO7OMtcAQNKNkk3Xag5hcLz7qfrQe
OYHABSKcjf7OTnyztVAsJL91tSlBuT/YvTEIGDkHxPAFQkyrkpXSs7g9yMOhURasgkKfx/cECDzw
pcW9wO2BS1GgrmgfH9o5w1a9Zu8v5/BgfBMcfIEsBD4KVoQJTi/CxOmm/WxaK45U5zjrclDaibec
f+rq8cbXsJ0HxSDSQmW8WJIYXwbCvafa0nfzjsejfKTl3kCg/jCvbxHlIvtSnAlM1wRh8ATFdgol
Q41kD+Rd+pIrr2Owu8lMm0IUW4QVZcFtAXUOs2zhOGF3CveBIli3OkLl49qgw9i5Z6KMgSk0FmNB
/i7VBsfvxzX77Re0f1CNLk9HEN3a1PZO3hTO5WU3nPRaKHK2UHRufItUFI/SxfG8nO15fHaHpO3k
WuvBOwT7Nnin+8sZy/JRe+QsUX9GvCc40tu9si8A+HyWvsXn92azgoUJrl5T7VVl8ge/n7qlgQH+
dXSesWDoMPpG35PGuy7mp/yN0YTVvQa8gnZq9CTqbpPFmMcK4GWA182+FSWXLZD1Nn5mTiIUwGwH
xBRtCIlnHBPxtxmDDZ316KTpljakrY5+zRvlUF5ViIdK006RRlp4gXlri+y6aCE3lFIGg+OfEgZZ
uAqr5Eqa4T8xIaIVwrT7GF+EKb5bMv5EaCH77rOLylQsOf2X6tzTurX5C2EwHiy2l4BBqz/39yKt
rAseN8jhC5QPnBevGmKiYP0jOANF8DzdCO+XVg68B6Lz7XsujEcHeBbxhR4UEiqnvZBI5OL2mXOa
WJkXV5WNvwR8RZnMlNprow4IrlDmVEoG+mm6YQWfVZW4Y8Bl+rV0gap5yOkVqOYt/VGJGKBGcdzI
NGlHhcqMtqNRxv22rchf3N/9TricQc9HnzdUOtVrjKDxEd06qCvHV8zKX+QJTwLHRpXEV2xdshs5
ta0Vw6hlamS7EJ/0YD0mSWigZ1qEwRWyGKwZ/7khW6BSlTfWrDsqA0MzmZ3UH4N+K3sROptZreuV
OM2Es1Goa/zuVInrU2JNMGSY2EDciepK5PZwdMTwElPCdM8E6b9NSBGweACYq6Z53ZuIcVBu4V2F
a51m5620rsVzAcDvLmr5aspIrrej+0te+aj3S3P1CaoQC7HJa0FryqmJh+HDpIOCSeebOizgILU0
iJdfP/XgtL/tY/q0nfYDmhglheiYypz1QG1QhVNohk6kzAeEOjPkwP6lYt5lkwDGS/VqwLTVVYxr
3vX5i2GVgwB6VpJDONwJe8WSuqH/e9lcLZ6UbI45xPITdmu1ITRfM1NQAibRwJboOQp73sBbIcUN
r5ifUCpe7zMIxWmxuXeHnvi+nUSK9gmQnDF4+akuUPjoELJp0g0EniUGjXTdi1LvPNDsaMZkD6qY
22en99ibhNyke1arpWWwHj1Sj6ILSyCGWLIy2Bp59xqWCFwmd/OCvrWxrYskf/K1grxQhX6tQ+55
oqts8+uSzHFG7L9iz6mBHraYPZABrLNjmNsS7XhtcTPtKvW4raYRi6Z8pUPxfWeuD8moZm/7Lxxq
ti9D/qzUjt/f5kk0E7dCbWymm5DQ/jEwIUNuXEmZPVZg5YqAGtTIYkjj4YMj8SealYHHYCSwXCw1
WoUFKdMFjJoNFkwSQtT0MN9oG8ZwEO4tT91TXaCq3ENOzJOYXnKzPKSO4OTCe9B6zEkBJ8dkT5nL
Nfw6JU5Z5VY40Eu+H3QYraHT4uSxIv3ho0gDNZfTLBfEknQIXu2YW3RuUCg3+gxGXy1J89DeWO8K
2Zk1lTJ0IFmAFHFDPaAUYfMPWlikxZ9uGrqx627IUWTrqW5A+AfMfeqSmx1lEOZMviUQcqpH5FmJ
BUC5hoHQdJd2wFtbdTG5Bbn+Bponmo6GWo0vDiNUF6CnqiNA2mLZiPFVoeZWpFFWeC1qRqgXCkv9
uevKw/TpaomgEzAG4aUUhoP8Y0tW2Ql8jrB97NbhsSwa84ezsWNDHtbiSZlzhV2CCIiSd4NwCkWI
H6FUHzgD+Ht+HpEeMbb+JZmz2iO/clP3rGbfyu9AQmYcLaHbLugLBEd+ESdosHXoz+sQsVMTE740
7SBr9+iJGAh95xO/pH7HDiR4yuGwLH2xsSE9XF4R5VZ0ce8h5zOp+fAgt+3VWAWLlH6qPG/dSMPB
Jt0D0bQnIL04t7VrWdp+b12yDrPwNMLkCq3O9r55hx/IOWLqrQewxm5zqb7KqWdTeAAey9ij9XkV
s29zi8ycPnIwsePcb/rf4glXtDZ8izRttr5bgP1Dq2cu7xI2f176BMtncCclIHRWJG0T958zsQz7
qoznISb3cgI53mfVpPEdGaHKHd2c2RywQvnvISGzGaJi0X50oDFsGnSCCtXlM3g5G1+RQoPXn8Qx
vMKQoZTArdO59DuO8gCKOphHGC2td7zQ2uEsjoEOMgwHqFNNQHJxJ6XnUZ1VZY8sRGxaIMuHhuTZ
GsZKBatog1qMyyYxuqKfEBHvxEx/rAq3vo1CHWtrnE4EQFgBX772lmxnlEXy5U7N88iWXD+DCPnw
MbIm8zAi83QRKKgIehgvBHwOttvrh+HVA52Xfbb3QyXZWm2uDTfNexBjc/JXq41qO80B/bnJC1rg
ekCBclkWeRIP/9c9mglMLT7WljHJ3YDMkmYCaevhqsS1bkMpyIyWcOwYZnZrzsZDft6Ivnn9lZ1M
EGtUnIyASAeMUtNQaUU3iWGReuj4JMK7/1KmoWRa/3ePKZfR5FwY66ZSayibE+mbroxUocFqHLE/
luW1vcdBwaKrv7aLXKi60PQG1fVRrFlVJfJwZdWaWD874M88wPRA409KIkyL84/2iM/inglzYrbK
+1wgngrPDdv6CJUO4LGFVe+3tQM4CNTpu8FYVkZQKLizDIeAVTkxSOXtiJQEPCC+1k7b3rfLn907
8DAllNULGvRvY1VNV5MmyxX55CYPBahAMghmHVqzikJKj6bslzG4ZEONvoNRrUKGBwbeZ4+oXbUq
yV3CZJSY5b4S8z9qmvLinU4WNJY2f/toYBFFtCuEFXr5pddsobuz3Ws7otET2QzNCh8hWz4oEytD
1wGBwQBiJKcGz0lN3uWrUfZGdfIBt0a9CwS9RCzGht3RTis/aqn0YWF0ppgSbDJpuVERBP9glyUb
gPEFRjUCQyMODRbP4pny2e+dFBnhlaiI11k5AtQcVoc/Wm0Eks1rYmizWy3H9E3ZR+5PrO2apsEb
p7tT0xAG5rLw/slmhDJtDHVXlwx/TfBpcfhUAbow/QG9FQUrbCQVNsBrGZhc6J5waxUqBLNmd24F
oDulxX9pQnj30EZueKtFxI+J6a4EiloZ0L6YKWStZJ5sGlP0OdReo27ZximanZOkfvEmvodrQ7aR
ZXYuYtrQriEKr+vrnJC4TjMznVu4FhB0w1ZXBbG/0FSRYvE9brT8M27/81cFq3xcSHprgtgqOrnI
xlAvR7Qmi3HTCM0sD7GParon22qwccgBEJIWzTnhQ051dDNptoqN8zcl5uAeVOe89/IK2Quyjw/E
d/ng/WysNgAZ7MIBT3ECHZ/vMrnDaKg6niXOCouv6HZRyI0zXkAFWf3HdnTYDSoPc9S5/25bG0ub
Mh3JUAUAbSryAVMjsB6UrGUxsepXXn+qbDMpQNBNV3/ke7KEghuNjbnEw212Hpc8JD8kk2iybczo
ar9EBT5NJfCCdZKkD6nXRYjztbmGTaueV/Etw8DjwVOK+F0HHNbf35KkEOVEFHRoJPzTzUDT0dRa
EZvRFxy34JB1WD8iyfpEW03pO0Ul2JxNgoxFb9qfzNn3SrgvtQKd4841WCp/ER3bnQqzZbWfWBY6
jJEyoXEtzb7cMruCVM12tbU/evi1J2dX2W7fX+rrB860TMm9xowBxtRNP7hvhz6c3YsMvqapSDV9
6kV3YlTYfUImDeamm5O8hQk08gRqYa5oRUclOjSKM4tanyO7x2cc1DNoVkfOod8rnOEtjlad2Pjl
Km7DWR8JQHmgpJ2IQXZx+97Q6MWEUm3xJXB1Owt/OhzOuQpL3DSPYUSVa8zfovjrxy5OZ0kW85Sf
wpR7mbmmTZPMwdHcDQ7ulfV9B4nd2MioE+wceHrM/VyhuNSlnzQJzTDCxoq/WoXV9XGtJ3HxiWmn
dR46up4UAvT1nrYZSb9L7wOaa++tqa9aKVkBRSXZisVVHvhso+qlWXtFwP/ejmAXN3BSpm0O3f1s
qRn1WyEP5k8H+GB5fvPmwUtawWhHD7JLktxOPz3s8S/c4hq8kpsSNoswgCo08SxUJNsLMHzJMBiJ
oOsUEDETQzXqpPJAh9J2gvXEj4iS+CySAvojRnMMB6xF3eb/QE/H8NwoH5lt/+TXWFxjs03ugoQf
sEeJ6ABsBBi74wJUzkPFUXLJrLt8WEJB4qV4l+zqWSTRa0FZZ2Ql/cxeQ31mJx0ZYcHMvKzpVy0g
WXU69OMmZ7SbgViVt07pGSZfcMgWmrr7ofg4K77AsywrpvQK+4Jzq0Cq2tgTiShkqsUjC/EqRljw
LtqdNuqd3wyJxp2k2IwnSDIXfoglmsTmxBHd0DIKRJaoUBbwINQehEidkE8eT05TY5sRVI9NKjvk
jkXf+1cZwyszY5SiQ9lV0z75lRCa0lkBOzeMbcxlrEovWbUO2BiQp+PvlXypGrrUdNdLfgiKLIg3
YiJ+LRZcP2xCJzbAvn6myaXhB0MHPw9EKHq9Rf6CdZT+e7KEvpabNb5Nt70DFUP7gRWCwhoo1LyD
hGCODB8NL4ealILPGHEy0eldzfgozN7Mh/qrWBZdZYcxr+iji0u26tG4p+WhUlyRBfsL+cXdF9Il
czOWyFsdeW825U2lbOhLXPChKv60tAy2nBvz3yACcSH2LwN9g5ewhBn3J8p4apSHtoT1a7nkhnFu
aUsJizIWvYPOs53LeVR2xQErfss0r+FEWTq8mqfcg7s+M2BnQBKs2jf1uyq0MYZItPLTmz/LusV8
0s8BZCUiz9buEkC30gJ2YQCk1imoKAqSFuJ78ABSCoUfHhmXR/hR1gYDQECNMQm7hm5QDJIH99v6
v77rN8tQce9M3i1Ya7FLxjhN0+Po3l1L2iImTf3J+OXBNhh2vSz6Oc/1V1iNcP301n3nwC/ep4ah
xzPCypvEnxgjo+VWyRz913d1xNg/lwJBHRdG/OtdQ73gGCeqJEOJsWdf6pHDyHtr0wYiXzxMZOZH
s18TAqP1CBherzeTui1XArSuQKYhUfymREn3ZyumED2OCkg/m3LOnblSQNu4KXR356E3AAA21fa+
xVVC0LA31eyZN0vUwq/ylJrZrHcL702DL0LdRizVx5kSz3zaUqAB7X571bQdUCKzCdUYHSCif9Or
9MsOYugXtM8Ds8yTaQGp4dRQ7JZUFO4fxXcR0q30ccgXIDuwBltFoQS6GwlH94Sfxf89sHFRlPTr
ovd6EwiAqC3V8L+ljsRp0msULFfpCmg7YWKcftAESHGlEKa0+v8iUTDjaHC3fVtdoN6OBPIRAhrj
1vmjZamlK0Rg0RbNjCY7F/PUksihgVK47Nl9YhWFTUZAZuLx9+v8iSgkIOmks/2hb5DUUIca6lP5
32DmzVoXkRA9T38Ev7A3yrXKi4Rp9hSXdbv4REZ/061FIYNvexFNeS1/1e2KMynJojGLxLZEayJU
f1SrGv8oLYQZNhvGRCCj6gjDcImFpFVJlgdfKPz6HmyhILlbBRx6SU/0FQ9Pn8QPqjly6jBiBtKc
3Pn0xpMQ2W5zmy5jbBkLbEysq8fXdy7adBZUcUsK3CsCtqFjoenUIy9Bw1l0qf5S3orsV7UMQaCi
EbKTR8Lm6T9JjKN+GlWBHcJ3Tg2QKu+SEIFuN79D2xRJASd2ohex3Oy+aXUGelMlsnYaduBv+kMd
0YpIz2jb4gJWg3atKL1/zYWnHFjG4AHkWIP0/oeno9g99ChhGStWZgKRyg7RRQ8ZyzlY0eNlvVp6
sw9T5JkU6ZomuyuWF0HF80JOvI4SQ+0N44etJedQsvFfeKsOlX/9Iv5hqWgopgUIVG1/YGS7dUuB
LWZmzbDoFY/F/oPoSVNvIIDtAavt0XTrg3M4HMGT4F7mp3gi01h7Uqj86ToX8KdWqbGHQw4uYnxl
NxM/ZuK0ScpW8Lb5PtFcmQHKZI5OvUbz1IJyE9ZA6hiEntxYeDFPluwnh2FVp+cD6Fw+yVj4Sk6U
B1E/AF/irAYXowesR36+UYk3eQyWWibYKd/2fPfiQFH+FtAELmO9Zi7O8nDQxm2IxvLPwPvnATKe
Rz0opfrAXzwjyxij+gA2GXT6Dlfy81RBZm9OwV/x1pVt+BWUXKvialQsjbr1p1jWTSA9aoXs4Bkj
lNVBK05arP7+1oYZQ/lCnTGQBrZ4c3vEQdeW2/x9ObIexG/BCo0i+fkx6Q9CkL789PaxkATG+xrf
USfhsiRUA8/VEyAhfmPRLLQFZblggrADGxUhk2dBRZmfHV3LMSIHocqoo/8f3taeOwyHlS3yndEr
hIzgzX6GC9utg7s7k8bdNRt/mfwH6NxB6zt4MMaFVgLfPt0olmFKqUpfAVllNJANEePRbxUCbcC8
9GgkRXeKFbpsU4/4nosGSLeckqiaOrDkEfPbDp4I3Bzu0YnrDuHW/3VfONRu+EcFVMG3tsDvul6p
qqOf/y7IT0QKPAQt397HpXMNyPkrKqSRyt9wxlXlNsT79AKGkyv/npuP9mBqwwj6uuArTqpi1TU+
vLh5cD+b/cJW8hC27itKhsD/pD5R8xYo6URablNqgRkn6J14/zz6DB3ngsUWkNXjnaITXFUWuLrH
olDi2xEf17x9/leLLEb9WA3ilj2/0rTIqxYwX6576Zc7kB7qBa+kowpQH51btF084ozJdmgckR8+
dxA3WFXxfYXUT2w9cQrjVdaUyHkRn30amxcv5A30QWNbKbsUeXAar1nWysYBjFJB2n31RGMTvnJf
yB5SmqvaK7mwHvGvePp0hAQ2+vBGCn4CngkKMoeqkAkBmZJkX59A5HWQsfx+v1Z2mqE2aXsIMWo8
phUZ7nAyqzJhaEBHCONbHLV5gCce963/0UDHvgN6toMP9ox0z61SDvBnA+WuTZ0RhoxauZL5uSyQ
UQB6DDXG5MIwyJUWD2eyfXTC4RVZOvQNWaExALqn/SU3FZC/8Cf0myVcLxIcsopMT/L7DiVy1NYr
FYjGdNO5cwdQgmBpQOumGZn5OmfdBsFsOvvhq9JrfcZm4rpQOFqi8P6Fo5GvfHyRLuXGM/82+/Ot
k5W+HkPp5Dq778QJVv8SIjrAFIPdDJCEwbTKOd6xKupk/M4Z+xUyWcOJV2/AkQxP4oghBoLRBb/4
cZRFYQQSSFblNW1HsVKOcu20nVRpzoZUO5Hm9eb3N85DeF2TB76BLUtS3nsZEcWeFjq9x7qQ3MSW
Pxl99vImSy74CVqoocIReKmf9MEnNAQzgf0l8DDP/Uf3ajM9lCppDi/hloZTJaHZJ/lMrqXA35xo
4vRu2UgAnCKf2gnTTfj4EtHwFiJB4zLt7htdTFewm/FH+NI9S1fdlr5yu7vwFHyBaRdo4gCvPPl2
9agoJwxSNMbkriNayjO64NEwwdVGjcVWbrbPY3RuaSAEGb60qBzdWVouRd/vXkOrBeh1HeBamVID
KQxXWRSsWDGDVTX2w66E693KTTyuv7OYj2LkwcWEYxNqihLfa8OrtziiJ4exf1k3Hxj6FXvog6E8
H3lAj111ObhbmRCaIvpgciLOTqTDh53u2pZEeX8EbV2/c2nPKOsLVZ3mW8U0U0NRzlq0crCbMoFF
Ot9vcRknCKaZh+f3MiIVk/do/1rPnrzatGMdSzr8MAR81fg6jZRzGOafXZ/JR1suiBLH6bNuEBxD
Yt3ckvFNeWjbUCh4E8Bb/ruqkcdUENWgzRm/cb4CVYYmVA5utKeEBdGztH08cfI8KBGBwjFecOjf
Yce1tbJiZMJfjKOUCX6vUQ0Tdph+vCxSY9UDNQ0uF5Hr0U1pJYwH1p1TyDXkOCHVMdiboVeji/aW
xgkrcEBUe1QK2pLYk7p1X6MBcNqTICPw9VUa9aLS/dSynTrfq1akpFJf41lkdtsF3qf2Zy/BvMuL
+1U0K0Adq+JQaF0IUxKowXPg3Tf1pxzDaUkWZiWfmgJb141aq7gGQmF6mr02LVNinB0CPsxAgKPz
CUd6KWIFyY6aliEwFYmDcEJv+XLVQSlexxBGbA8JPBdQTlV9+oAgWaydYVryLcStXkJjf+K0w5eb
2BsHn8ac9DatyOTwegdWTXKo8Ibmu3PAgrS8LdVrtPcqe4iB/Tvswfx/bGBqFV+wiAdSxCjyyuAD
IqHfpZtzxY9Z4PUlZSJwgMZ3dWQJCFC8ABTmLvQvq4fICUaUHS277xsExv0WwYqKR/yH0xtxJ+je
V7BG4zO1Ad0k4LZTWwb0Oo1yqI4j9gczj/ufYdhCS9pI8MP6idc8JmITwAsdfzw7OuIczBWuFhwl
0Ly8iW1GtObyEfECYYZcGD7SOX5voRG9+W4jzwNwCqHYDx1L2CTo0PI+meSQ/OZI10EhF3yNDJi5
+bdTV37fRnO3WQn3XIko0zHFWkoZs/yJDJna4tio63OwS2gAlD8fhls6ZZuPbkJRklccSfV2/E97
0DGAV9HA1nPh1LCP4IJPh7AGD4oujoX3uYAM9uEWNtX2EIRMp9Bi677WxIQHv7D8CWESPnYsMYVX
wu783PnZH+yugPCGo+OrcfTAsj0eQRlzzX3C+uow7RltLEENdv8deSLCNSsW++rZByL16fvvSJiP
6c0sabdMlDiCnK57wGj7LQBRTZiZxxQsTH0HWDnH96aaZYlT3DpFbdTV+vhaj/iC0KTgU3LisEIu
E/QAQIGFhvaOIoqMGg9C3FBbJiagm/N2OEQTCi6CR5NANIy/jj72IqQ91sUOawnDhgE8Y43Lcjao
gov2k5b9VKJS2ZyZDsjafUvQupWDaENFIPx7OxUZv4lrg4nNoVj+SZ4RWlsbVcAjmZv6OwEUNQpI
Zzm+jJoMPQmUeIT4IcRGdN4Hc8BfDvp0Pu54J+u3e3CY/yFNjcsA4iiNSE8h5FAscpYJa0ymeHAf
8U3uZ+IF71uB7Uh9g766KOtHdx42vFHflU4uPSpqKPI0rAuDNvcnntuifKPyIWeVqA+xnuF+K4fO
6KDBuJudbjaduOiQV6sR+/944N/Y3bRtduuscFCIHXsSUC7f6yyaBfFAXusZiEdwbgEHhErdmjPv
XY1FMry1BnDCWo3aN4qhFrZ0Yw2edzPCkf1fTrEehUBThvrWSZbttdYSvZPX66lrlBx7KoNXNEgY
KT5/Nw3RMFfGyGOAkQ+x5l5f5xsdBRJjFo7ywfaBFaA+Gk2uN1L4c7e51z46ulyMhBhpjPZeD3T+
cyWgE6VgSCaThgdXYQtkQGGj1WWaFUe774fXYveIZRbFGUQhZP1py5tIxAEzI2lzQt7/bgXNbKOa
eQ+vdhuQsGDlIQxb5JDZjcGSpMvS2rucKvhZsNjHYTM+i0xWW9CDqbkXE2d+N/DTCH1YPmO2Vnmx
rEivBPxRtWNsM6NsYUMH3jHh7QIJFNUWacH/VCVGUPx4vDJy8MQIcMZH/4PjwOb2yUomFWIX2YKo
JA9zqYPdEImToxTplBCOSSOMozZ1avHcmLHgqtJNXGKA8GoStR9zEra2mdRhulhOzXyIL1CBTTHf
PYfwjevoNbNv9IBt+Co1UZ58z/d6jC9WIE4XNrs0/igBtgHXZfhPXQZWrcCRbH8tRrHpLGOqCJn1
OrydIl3y1cVbF6sQtvT0orctzkXafDdzHOeRB+08YzAYrzAiQyqMjXAXae8HLvZJ3i+LJhBh2adM
ki4F4tjlRQ+kcafuS0IRQjNaGoCtGjEqyOiNJt/ponoDGpDU6zO+7to3H3u62+CF6KnyJx0i4pWO
cApLrlEou7onAVD4Zhs4yapz6P9GIS/60pBnA8tfWHYiJFg40Vl4+nx4rUGmCcHQLeA+FXnqTnHz
cSvu+pHiSDfp+pi13sRINj3Sf+Ny798PgJILmgLmGn5q08w49MTdVDhiN5wQIT4Ji+dl5ieAH1uZ
Z44Hq8qwVQtiM22OvmElJqtgtMBlGCNq2364VlIavrwLUvbnesOxKAvrxaATaTpEY5LjK4NI35Dw
zJ81XHwauyVuS9dbImBfU2ex6xtjR8JD4ZaMBLcQg5fM8tZSoSnf85aYRalir58y5RP2vGTHsGiO
xFdIBrjXGlshvYoUe9h4IK9H7nYvx1sisdv8AzaJwvx2WJEwbGEMzyLlaLttES6ICKK7MVjN73Pc
/yO5aIMEeSYM7rmn/1MRRkHad9DEkZRJR0jzZMOK6sgyjuRac9RMKTTSXuMQxl4mcJm6N50srjAl
Ft3B+fe5rby0PeLMhWJLNVwUHUXSAQpZoNDmIN/9JqWFPHXkwfqyOoQxg2IqJ8ZgYv2PZQW6wbO5
85nSOKX4+wp6E43piBrYfj55TuK/2YB/t0aGIYukGimnm4wbwdd4IYuMzVWJlhHtw9mQ2MzShSxA
vCGPlLSPqUbjI7z2dUV44MogBUm2RnxqhzdzudzUJ5gvmEhtY+SFeSJzJyDCCiet7dYbGjfwhqwx
YYu+caGLQt+/H4I0y6+GOirz2R+dlOA9WkN5v4B+rE4z66o6w9nQtnQQv1c8Sb6F18DkjI4VsoZb
WlyVlpl7xxJ1Nk5o4MioNQypVU2Lafk3jMEvgmDmxz/rc7aL/bDOewIKdu8BMNXpqODeW+7D++ja
HwFUMX9jeQsYQ7ZShk9ePpdb62SUrF8TWY4lzK4GD0NVuOFhxqeYVFKrQQ8Em73C2U937En6/eUw
BZBnAKjuJGDiWukN4NYwGXs2DM+1BKl/jP2dbKF4t1DjBGzS8rvX/yWqzpV9DIUoJSrPdzX2U77V
t+iqwUoQhILe8C+gR/73whdYnXaHnrVwQpCAg/G8SX3nv7XaLsZhuG4n3umk/tfjgmI2uKH3ckKm
C4LhsSwRwjUXhyPwqBOexPqVOKdybCsKtezNUnlLRoFIR2Av812e29g0w5hn7jHNe6Dzl1UhLRRk
IYqZnYMdhJ+YY7dGwTiReEDfDUiNtACXqNM6qeBI+J7kqTRmP8FZnJ/rva9xI81sEat4no6TdaWL
tnuUssM/+DOYunpjXpqOFmsmP99EKKYITaetZVWDYFEldL1zVZnzmy0uB5oWGfFpv4pcwyAz5BU4
3UraANSP9rlDXUTsremLDQl7LfEAY6+rk4MRjuajHRsgnfuGSr+p37iDthlIXEo2QBhNZlxHBqxb
ADOcVMoq9ABtdhUxXL+a8EMbMqjaWp/VkUaHveUgCi94brSrwji9zYHMSMJOTL99ZdQsul8aohpL
gTbxpG3qe4R/0yXJp1xjTxTT8CTujFS0xoNSeFz7wqsKWpM4LmiQpmy/vhNH7FvvPq3n/YXS771x
/2wqMnu+72sT5K2UJkEwWXx+rKYpN0krmh/HSBOC1CzUFYAFmJgiQhXou+/XKy9wvUmDqBMD0DYs
sz9r4xGZEcAKGuEygKgt5CKV7rc+TAl2a/YoSe33MC8QK1L47avXWcNYp5/K1qDGFBinEH7W32xC
loG/T2SEomPxmyfmNhfY5Y58vOS43YoEV/BvbytvxHKhigvJKT5AhP1VtRrKNMLbClXACsUnUU28
eNlHVe0wgj4c9A25JYAJeXFC5LDjNquEHb6kfj8TO67ZAjwIKlC0kZ4n9Kkjea8eJWMHhofgPjbz
b2hrtV2i80Anfo8sLkBBcA9FVPi03FYF98+AV9j0H56wnm24xiBPIgmRttQZclZt0CqI8g+m8m/7
JKLPfYzSLDmgGegATWEL/0kER+ytBTcHVETCFaI37eOOH4sdly721/4kt+/25qQ0EJiJWTCbYpq9
2/YZpmYCJ+Eyjjy467ri8xiraiqD9j5DiB9bj0K334TdnOay1Jj8WqactOgCy52H7LQvg4g8uvoA
Vvlgw52aXm03Lh8fmMG2u9QVr/vL7ajXXsDnKYvcBRqiM50XI8T5qTdB61T4fIsEtV0/bcuPEZ+r
BvKDkz+DNTdCpMofFGHwX0TTkX2C7+A33/RXzzxeGE8e9nnZMEA9k3WHQ4k1BhEqLVWxz2mlDLS3
io0eet2Cv2lBb5Po9WJdHuVxpJxIkBbmHSHyeQrH0ES6u9Ix3zINGjrkB8ntUnR268aR9AFWVcy3
VtKkldaDI391p+RV89r9LCnKmBDGXO3UlwddjN2ZI092YmE/cPraffn2ZuWlvg3ktMJAKCJzd+ZI
nDKGjwn1fhuscJFEsdnZZiHZT9RRAZa+MDNfNQDghJeLdlX+GNS1mFV+RrbKNGn/QYaTWKLdZE83
4sDEkw2L3vjBg0Km4/eD0nJ8yytQQZlPA4rrj6MWSbJQvAXHSIRB/M4RQS1z40wBjRN0bbKKWB5Z
oj+xMuYmCDDLFCuKnscc3qvLzGDjetWjinHdrMF0vhFV/Gd5GgZm2BTb3omXFGhumYHNNpU7PrWz
DnZEsobGkYWGSP9+dZPikCthqbqfN7Eum6y4S87KtKtiKIYxlBAnD+wcJ/lVFFdJGgwhovkGB+Oh
38ilvUdub2ANUDD4PQefuoAZEVE+6ztlBA8v24ZssU32MaG0UBWqwKzMOK4eyC1CdgXXMHLe6Thu
Y0s0K2He8GCmYc8DXNsmShNKfNoh/Um6LYerfpcZJEQVXqtfjN8iZ8NGWbp1aDCrVLmJrCctmW53
qhyjMUJXmq2QHcQJxk52bkKa09kZYxkKN6F1sa5YegOhTweVfSa7DQmMfwNCgmdGheFFR38rT2U+
burU+Dp4dBQ8dva7fH2b+Uca6rM0Sz6QN+rl8PnPAUrn06za8W8ucR5o4TS5HuSHl0fy7DeMV9HM
o8Vn2zx0k0MQLEEO9eFZ/w10ew5qE6B3uBaFEFPsAXTrbm+JLKGXWtocC/F4WjkAeuDwAh42Fj2R
gSIIyRBbA/3vGMIOaroGmHGxJejj3JS0EqGskrV/OYlH9iLgRUwpJUE+mFw31RIM7MSG5lj9veIs
1bWPB0Xt6yutNPaJk5+DuXL119V/93r+ORpYY9EwSBl6paw01JK8cd8EYb/t6pd/n171t6mpeRaV
/yK6A5l9+laL+R70x2YHnloT6Ff9KWYD2/Q+VevwKWvGWIszVN3K7/Dz2sh53LdOCbinaLskES91
pQkjBITVR7ITvp3ffE0unfowpA7GgUg8WlPfOTmaGpvkk9GOsiw4madn4ko1b7AjtmmjoDMLsGbt
blDWZOCo8UU2r3PXBdacUU1Fl3p+FZ+JFtqv2bzmwQnqRiwzBnZGBOa/kiLPRfDC+iMsFDAWlmld
ZAhGV5dXY2ejgJmBOaAZmEXpx+utu6bFnzfwFhXlb6D0Dc3HVf12gCAuffrt8znCyteQpm0QRQ2L
fZDd0QTlRznUQZG4JRX4WopTsPgTE6PLBA7tIC/XoRquayDZFb/QyfGUHgh0eqD1tu4j+Cvzbgcc
E579KfJBuq7RO5Q1Zx0KhZ8WtpLolkz8ACrQaZpgzQ3MhgiszDpcdd8f6oVJN/XhHuqOe+ajQk0c
r75YYkVoE6p5WVPx7o3ZR0EfsiIKQWi65gcw6lrPxvw5OyxvoWaQ0abZk1Mqlu9O0eUgE4eY13yz
uFKfqbGGJUhPZx30GcJ6fEi1oiRdk0YKnfUnJ7+jnL7dUO4gX8DDtTvm5oc89W/oOnTPdFoILS37
apjrBkYblqtlegr5d9zX3nS1vKxlkqXSb/oqB4vAf91LysgBzgvM6VnyokwKe4hpySkvUhGt8L0M
QzeePND+94/Y0OGnbvN5WhqLiEqgaABq9V6+QrLmKKUie3C+ZIHqEh39FbgXkRDf6iRZw/l3ftFS
QT2la+nqmz1RwUJLIpSHaI+8pg1gL/sos7tVJISTyMiXT32kqfiTgLkrBudRxDPZkXyYVwr1tGRo
oZO6vfvKvzlk3PIxRJ9f+gEJC9Vqbq7s9hjH9L2NVXSXkjkoAIo0Sm2kdUApagQ7I63SWRMyWSku
LofDWASa+Ff2maKatMzHQdANH/wuEtY2T+EQdGAgXdnw3c4EGIkcN/yiDrNNqWvEsVkUekY+OwHr
RJ5Qz7xwNRzpWx/Wyt6SkhdcmLIDShbHgkTLyDxq2r7h8bEEEMNhA64HUMzbdYzuCKdHPXJDmo3k
SyC47KaAJNCVTfOn0IpAtrgODpcH6uD7wFd9LqizDBluQvpDQdIjqoDO20YX/izrUQytnYDtPHBf
D+dgJVpJOmdEqCZZ8hQWNLsQ10odGp9q8K5xBbHSXOlyhE9UUxb3ZnKiRn97/lbSwGgTIzrAvYt5
hzLp7ceJETLYauyADtIKVrwM8rw3YOj0E+ojut0G0NS3sSypaIHLEpyaI8JM1nmLqnGV1FiHgA2l
aOmMm7NPLYs8f+CD8aj/KgvvVqthgym+jyPOH3dMkbzdsiJqQEFgH5FriBWfS5wVhyrGuMv+vqiH
z1fh8PePlHIoMnafqKo+ezSYGBfzFEZSzLLLkJADoQN35+xzAzwemHu+OoiX2Q2NxTB/+V+vAy7o
3fQYX1+joQWbFfA/+mpk4qoOGcsbX0dFF/xkjyGaP2OUPVVbD3+fRY0TWercOmVvWNOVhN/4Y0FS
EENJfVugb6M+IpqPUEZntnWJqjik5NHow+AE3u+pQW73Qm/NTsWBq3r0Ti56rfKGpFzrEkEtRGXJ
AJcvjk37svWvGGrvs+hEf3ysYlAsKWnzlhJcGxnNNEwNZlyyj4s/KK6Wxp78H4sOEhxUlvbE/kaA
spsNEu6zWU6ISMhZSlmqBZmCXHLDz1kUvx2jE79rJHK3p0ZVK9zII3efOHuDRVBG0JnmQT8YW2GD
TmDcdxDLpvPkMbM38/w10OH8wUjjaWt1xpdqAgdA6wh4mr+ePWlUASF95RsSTvUAhb6BDafRNrRO
ltOZaSWPERPi76SDaAAjCDvI09dqtBDOUilZXQcdNNHBHUQKlrbuzTgptqQiIQYnpe8PtzAc/LS3
CY6Em31w/lSulYjhP7i4n7cdk7EeYkAVTOx5DA91SfBLfIGEjFpbgTByPqAGLrQlPpa/mSpxPndf
flBHskFb7KQYt7UMx/Di0h75JX4Nwhmf6Pc5zmQizWxRNnzppi31xS+8rmU/lIaZ7JZvl2E/FU3V
yspAJdNLNoXeEzu5jGlPiQMw/6d73tTGb+LxyJca+I30tV6qOgJ+h/iAbgCwOjEs1koVAHVjaFEZ
YVuqwAe/VeCnPi76SK+K3AicPRTj8PZZbe+sziYHS5A5ISe177ASP2rWc3sAlOkd8jBshaJcSB6P
SZ0m7LKeeDfaYv14ZUPLVmnrD+qmrp+1CJ/7dm694Uk1EC8x6W5GiEQ7jT2/Avd3j7Ili11PDKPV
FcXhqzHtRgr+SUFEsUzLMb/aBHFO1oBZfiHVxXvlchCmy7sZpilrvemkUj1pbOxlZxMKkGesIQED
I6+9zjrLAljzqZgGZ+ZDqeh3oH4dBGz7K23BVuKIkKpBCIlQQKp6KNZ+kZQlcMGQhZzbja3dk8li
0WmHzq0Nyrsv5vplt6pexiBfge7iBi286pN4UIsqxqlJ7+msvVz/j+UEsh6SsFpOddbhsO8ml0+X
F8NIrNXRfLdxJ5FCt9VgiUjfHGxBXDGRoY17MxhlobMVGE9sF+IviPB2W3oN+Yn0hVTnhq1OOIOn
nTa8MVaeoT3UepSo4y3E/PRFFeAAgB+xMqJFt/R6dwdVsIlj66pNZAc+P6lxjxP31Fc8+vdHvaPl
fgaFH8AVpa2j624EbbMNIe+GRp1nhmRcMDEYwNRdNTC8xjMKMdp08IH8+QTxAk9scUxr9XXFDTnd
eg4ckUIkIMCRT5JV+ADuJ9Cak9sk70lTMWfqCQnlh67UtIvaPtcXwe9+5IV9NwiyG2IMe7m0bzWE
UTmskUJ0F3TLab7KH2qsKb9c1a5nKCbLOzZ8n8zSsV/aqgsl2VtbdrCnw8H6xGqbc+FPxVukNYGy
opOwh6zt6Oc0LKuCA8V3myhaOfmmoZijDejc/Sbqab4c6KcmWuo2G2nVoBCzNJfmDb3INSA13Mfn
2lHDpqKU4cfgRR93ldGESqGzC8x+/Wrr7MvAKmiFQWIey9jR7tdp6XeCPC6L13FlbJOhUIkYRzg3
XOEiWSOmXAtHtf1bf8P6mSlQvgZRd6f0MAbD9hnOqGFgfg7NqJQvGSGQb6HXR/I6zFElsKxIipYj
Gctuy/b75Q3UQQBMfuZ4eh/qqnkdnzU08cDV6pDOOKCke3zGNN/ZEvhoqAWYf8XICPTmdCJFbgL7
G+ZU2jx6pHxCECEc0EuPt7Jn2SZHV2KxODZfRTBRJLW1eYE90drN29y2Z8xXC/RwtLaFAqyzDBbD
OU3OcP1a6uisAmY/cDi6hecdc5wD/qOXZec3QQ0vCkyuUpiZmysgfDfHONJ2qoCGTGjKOhmelmRb
77drBLUGB00vGROC+QsKGdMjGYrAENbYadNsBqgPnpzqU7icdXBvQbgzHd3AoBfhu+jpSw6acCWT
enr71SYF+SdougIwu0qug4reivroo0fKfSSW/AZfxsBrXNAoxW1qZGKmD3rUFqqu5SSdoZ4j7gog
0+74aWGJzvl4AREDSJbFCb8GD4m/AfVpbndp1SA0tu/UUG3Yl79fiv5ea0VWOjDUD79pzjh3mtB5
5ikXi7UmrZaOStLrFQp3HoW5xOMTx0PaAS4ZMkwqBk7GWoQlhloEASDBhaX/wxHSSoz7CzJzNvIb
K0KhQqQghaLk2CbARvctdMK2GIO44SJwxvitD379k4J6Lw4Bghv/6K0ax1puIiGHiPIxKXCozDnU
tx2IIhnnMTQejaUyt9EsRSTN/+WPs+/Sxo34eYwmjeoWZLlEr5fQpG6o24W9sDFeJA1WaclFVZ4o
r8n3bIlkTYKh8H8VzAZzgENP7BumbRn4vmWj0GYpSX/S8BzLxiCLo4sbjHOox+i9rDFpoTepHrZD
pJQuEAY5EiPeP0r0EAobls7I491IB+5DeeJoC1YI7Ly2VkAh7W1xMZgUZ3QbGtADzSvgZQ6FHWu7
iK/gzZ2UHyGzsjNosMo3YV0gpYtUjKnOqSBXrk4VvEW/WrHJ25sTD5I24ROnD4qhv5oytiQivCR3
meQU+/vu9Q0tNj+aqEMJpRIdp23VMn33o2Jn0N48tKnxSRhSk8PUOXu30kuX1NwLhbLvPyPNw/Up
Sqq8tq/LSgNcnt3jxOZ26OyGmyuPWAWH5kjPb/nQBKeHnQb59qE3tzOFfkY9Ba7IsGfU1xFMxZ6o
KYqlvuTJW9nMgqZyG/XNTMqAFbHgvkdvpX+fK0u6chMB9E0VrRaZsNEIE/TdfBiff/DLU8dxtvE3
tyW+VykVjBwO5RxMc3SG7ZMF6Mf6bXT7ERGO9NFLskrXyTnTf+dHaohP7s6DAIyLLwi9ZDOUBZch
I5EetN4GAMb7ksPoe1N75ETELpeel3lFjSl3rZtn8Rh3bTmqILBXYJ0TBdSOEF8NKFxCHafePYMc
PmFZw1v4aUCjHu9df8PblLYVVQvxosvVE4r3fEN57zRi5RK+3sn053k+5e++tEEt04r/zXwKoFdo
gmslq7vA3a1OAODK5GdGhtOVZ4TDFOMLFW41uSlsSjKI9P0LPmEJFl50EoXVU32IzeP/y7y9tkwF
vCkNx2KLou8O6DbTTAaCDtmuY7z8qW0yugDfOtB3MSxBaw6CSPaUjK2acMy2ztcma28JdHDMhaHe
JtAsRURuXcTMV9xs842YKUlZ3AV9qRdZuBCF2uBN6DTE7VSMHIGy4cKXGcdDbQxUqq79ChcZ2c3C
Zo83Bd19SNl3nxwyAJ3UxvWU+tX9fMEIcB155+ieYuyH54pmvUax/zcYJ+5+I/n/duNwMuxSG9eX
OSP6CtT9wPl++wcv7UHbUcXUw2J57ag7k9fSg9zDM5rCK0SCFLdoA2+GdGiGTTkFFc3oELxJToWx
qP+9q3rvVlDcgTFPP5Oj4oj/lScrK9tFLqN6SkfZQuBf6xQii0IgMsWg+zSFF2s04IE2elLzFzKM
d47ehjR6uNYakNe4EnRkYjD2myhFe6xAP6Bz0CMNUasDfguJ6tY9wlvywLIxTY3XjFBmOYcg+KAi
d8exwgRwUHXBX1W77H6U1r0AH7icH32Hi4UwXPt8EPFvGt3FkXRyPEF6LlcjPbQJ+Ntj1CPoAI5v
DeoVa/2+n9j69GqX1eO3GxRVNxGzxy5xPSKmdRtk5oQE0+Htb4bCYNCtRpRJt09mJ2MRQPa51/AI
ojSxzbSavLkz2P2eLjv9k0SEuXhuq9FKa+D6XA3wZwHmcisIoabmWULuYwmwdTgj4sP62ekyjpk3
/suYYKjK5wA/dThnyFqv155HkYVjJmplCM9HttRPpfaSrbXzv2a7vibhoIm1Adn7ne4ECeAmeehQ
plW1dXgO8JUAI6sdrVhnalvppT2IxA8vupwiKV5nxLoyPK0IhC1YXzkXaNPzr8G9gqr5kIadSE8O
eUWYYqeUgz8TYrV3FmeJWErcVgX8hjvL+Q/ZMoHBe43WRGizS3AAThembRS480a3LUkukpGTQ9Dd
GjVgTdEmxjOvtiQU4sAr2eS4fi88y53MDmJZHqmzzyyIpIkdzOjjnMra1F3HRRUbeJXITDtHPpDO
r5btc8rh/ve31laiBoKzlhBBcrMJQ612GamwDrTniOCMexLnUxpcrWEGdH97Pw7ZUZWIy8zOBdxq
o0IzC9k8pItZ8AzdEkyT/zi96aMGqqJ769/kEkcUwqOXNkoNC3DDvLV88W8NUurC5fuR/2wsvZLb
YEx3iQd6pILMVaLNo1ctJSVsyz9ueDV77N0buCKbId1pJnt7qRuYDmBk5koINkcwQKO2R2zGEij7
UeiSmeI0RNJRxg6LsDK0RLBvyFqCe36ySuCs0rF6RaZGpm3QIk+wL+eZZnkKdN9zCPukcUWOFMS6
ukxHKfaGvwXNuN2rZhXTWAWOqXGo7u41ghfm0ZeCJrB5/ykYMc9HC/PMGzSpD0oKg81TkMCM7cTy
b0IzvR6gSDa29A//jFqNebMgVg/omaYPKV5ksxfpIpKnI7f+UBpWyfYGFVgE/3NFDmri0zlLkPGJ
41owdTRhF2nL1xGUeUssYNes4n5ING12yshQ1xkcKvQzuLOQkJCVSzvTTnSRaD8qUHYAJTOQsEoC
R02Zrvk5ORPYX5dhTDhqHJ/fHh1MfnRlnAaReS3pbLOFCcdSPt0NEtVXY1bEeMJ69e698ngl/UAM
T+NEHhkAzN3wEvl9eMcnngo00OFSnwBlG18Xpau332Uv8e01pRJoikwYQ86F0nL4fYrjymq3hhxB
sgc5oEvmafZcmH7ci0l32WP4fhujS9cWzya2r7r5WnfoF4bSgprvzpHlPoc5dafF3ARq8H9FoBpG
CkXvZswrxwKfXAWjSNfVR28tSMRHaGVghYpH83c8wUmBUTBJ/fjeZ7sz7kj4iS0042lNDdDNkWEw
GtkTACma+U0pQd5pVKRwOgFov0yvkNNRUganW8tgauVWhBKbzGMDRhYkHrAkgIDx6Sc+y3rB0c1S
1TOD1itzsNQHEkPgZiQMdMBx5Si8//OxbR0wfzvrtCvgdEEr0cZ+zTLVROp4iyxp9eShHdRfg7bG
J8YQv38R61JVNMteSqfUKo9FgnCRh5MUZBXRIzJLqpn2ZpKEuwwwhFE7pqFPfLCZxn9lAmaVHX2J
6Z+j0UG+MyUNr4dcIHaowluR+7T7Ec2MVnVXLc49zzoZDnVK66mNBA2D3bA5F6fgp6vS89/uZimW
sRxfEBZvOk5Sp9jOZ2uzsf0kl9GP12S/41U84u8mzSxqBXp7Da1w76tb63+OdyLy/JWwIUaWGW4F
N83VAAsob2VTzEDAi5v6TWt7iqvoxGa7qgz1mMpqyZElDEeZpGO78YembXQ8lFE7hzmpxzrCWU7c
GljxTie395jGJHmhkZhBbGX+bekTo+GTXCsv59Wb8M6uu6M8lnjg4t3EIDqfcfeO7jK+VYByAKO7
qmmLk8iwIjTGI77AqKpGpC8uexjMPIrajMnVIi/f1TsQDAsTpeYhoxQjFPv/AGfkoV4O4waNKYU0
MRExI0P7LkQHWzLRExP51cbdjqzWGoGwD6XHZ2UNvZcKViFHO0neLfuWI3WRUSZHYZkPJTUqT7Lf
HuFUUFWSfu7tF5EJdWoJSxymcAjzqONXjrazynAbXkYuoHq1vgjonDhF1QJE90qvLnB97g1ohCZ9
P7g9FSNM+TFwMrZEAcae0is2DkA1785vrttX2INLUt7uaW3nMzK/q0m2UmUA30VxK0KXLLn+Cvc8
3Kw93G/WSeLNw+Bvgkp3fF75gg7sPlp3qRfzOaQEPVwmoBpdbOpFqtc+dHjyzxPp/59lHUYC3puI
47WJBT0rJx9yHpzB3YgbFcwnqiiPFBn11lD2NcH7WQpt4fsBw4dxh40QHU0/uIE33VRqnY8n24FO
eE4bS0Gw88eprF8CmB8u5YR9W8eTTdX1S0CNMEC4lITmx/D3zZS/dMLRae5oIcy1DpBcbK6X0HXc
U3JHvV52oTE4U8Slpr6f1eRBnz3/E0i2HwjTQbH9zUF9S6NP86V9WAMa+25dM73hz7o8jxQ2N9Ln
hcZXTbjN3vdN9Slnr5JABKe9Lx6FAXNcA8zx7JWp6/QW/ly9b2u6Ox04hclmZaabekIfBPRDrssv
DWxnOkgpsMrrp+bidYqd2ahxe80SS3EcNxVl3OO/lUPUc1IxLgfwhnjDIIsRERpuZBAQ6vczh4v5
5GxDNL6NKqskgKML3glIg4llZFH57/c1RvSRuQWosvPXmhMduemXDaK89AOZW+tE8xHrRP93hZX0
jQuDDzxLib0+7G2BvFjsnciS/lAloeXHFTW6e6BzbJcwKbxTafDkWH6aqMFBv3Pene4BWmUPOvWm
jfIlfI5pZxpaIlJfqaJ5zfCrUJVlitdVqHV0qc5RC81R3Gr+vUY9cLlJHNU0te+3EUloVKsdbcb5
wqIz6gvPitYpdPyFlJLNpW5uG1VRfO8N4khkKrivqJdFY+A3qvjBoH9k7KY1yZ1f5ARQLiNX6t6h
xwuqQITFssKnaZmXmAnELObvv476tRMgQNw6UB3WAqeY4gyzKvCR5duk0nOGDIChXT4j+UHEl4bj
P4GeWFGfntv5BVWdjnt01XgVwuFYZkb849Q6WB94Ak3UOnknOOhMlnbHnvgHyHWwCLQ+/Wrow349
wyiQ+2lWB1YYVYu7fA10610KNzGypk813KlgxFugvYJe+trj8B/tUUGf1fh9VhlEkfraDpqP7eW4
tLTPEB+HvG1WGQ/SwIO0Ky5qWhU0vMq1oR5foPq9yBXDDnc6prh38V0fSsFkYKAXdUnfU6srAHw9
ZZaB+wQv2wWWARwZ6P5TUeLwa/se9uuaEBfPXqWrkc7dDoCdIeI7s/x+/g16AWyR6y8y81SOOd7g
51BJTlC4k3I0qvPa+pgjnOjRbhUWvb8gWjjDWTrnAKYU36StFIAGzMSqywMTIq2EpEY+DLt4nYep
5PGqmG80ecTkKKJOYXQdEJJ9ggDRsHQslEUjS64NLviYryH7swkTAfaPJV7hh+csR1UVw9Poln7K
CCBH+BhWZEmDpidMG0LzO2KQ3AWUhxN1QJ+rhX5UgLkYeV08u9Kef+T69wJ8B0I0iuzma0nIVhmC
ES7VhvKUvW2cqfaABiDi08iwSQqXSHshMFo08pYapgmQv/0Ui4KG4OIVpFsCkI28GBcZgFKwJfUt
i+Lu/K4beknv1PAp3Nykhsl5It0b0binnpN4ZJygrcB3ZOpVmmsAQ3bGVoojFEMjn5HTAmzW1l5b
suOL36X1meddaK/kGqqZAkjEtYvyi9spneC0CnWRKfYN04N85bHUSjxQC6X/f90lgSr7dgficZJj
HMRe3By1Vfts2XE8WtOtOyF4jVWmRT/D7+bSkS5anZxKqCZlw43HYOfPP8ooM/+UXBBu4nVJwP83
ml6ZeSZqcqf9z/yn8sGRd8Ep5WITSWwgFGs0B3WnVQsvoAy+lz3pb+pbQQex964CBVN89+0RcOLf
PtvyBI/ejL63dpb2gXjVJvMl20SZcdQjKm7qgV7tmCioysQSTSKDejHPoOBI7HeE9JR2WlNbCrR0
t3EzRHafG2krba5gOo7c32+BTA0L7zVddglie9b6aqvTHsc1n+RYdlg8lHIucJVCnFm+eQsDkloX
9QqC7zlfS6GIWneSmYhwAbwxJMcc0CHepn4u5K6Hi6DikbZyHm/GxKZBoig2fsYj46WBJmQWF61I
79fr9f9ncyHzHphw+K9Qamu5GwL5gdK3p8J+NkZWnkTqyY8cxf7kYi7K8GTjgDTwlMuyvu8y8DHR
/MfldiSwS3+H8nuklPKSHFFQav8Qf+s93rujUu4kmhsv1u0IabBQ2O6Lw65eKsC9IUDPe+s33JLZ
ipI/RAQpDi5QPqv1Q756++QhpC4iOjec5YvCB7VVEEH6OSRF1I3RdPw6Sc9KQrfDDBNFbJMJjBAl
FwY/TdeQeIn5HGIvuHFu0gtC9yIs/vz2mXqSM9Ijp0EQO8Oj5TSk2Csbk6zdQsCAhy8nU2Rhw7lZ
XvotO/jcEmCitKxtEJUbeD+0cVh3iRDEa9XJWAvsVHDQWMzpqHX+Yro3uSgvN8kZNRtEhqjkvZxg
zh91Wew/U/iSE1HYEL7am0xn63SrPkq4vcCdgNolCL63VGt0IYFH6uM5CqhhZZP4gh3vPmDsicxp
296xpd0JZGpa4PS+SQRNg4zkPSYWSJy2PxoMn3oxEoqGJxwtwlmeetDZdK184GMYwtgrjoqxtfvq
pYCX7RgZvXkbPaeMK4uw0N+WM+dk3UmFZdh02rsvKU7mhzIvzCG4f1PAk0eOGTMGH7kfi8MVW32B
e46mkWYy/RJ3Utz1ZmJ6JBo9Znzvud0r6qa0L2p7gJCYgvHpijPrCp73LBy4oWApG44AyAiHb6TM
sWURQh5wnIf6nU7dsMc7ia95g0HuZf760fUkRGQf3Hf7GiZD9p+1g8YAhCn/s3VKgbb5EzILY3RB
CDQGFunZEnt2kiEH8RvaU9gGOULlyGTYM0Xwbj8Wja6y2ZqcWOieN4psLVccyAoj/l0q6fWBZiv3
qMUe3MRX34VgHP+iuSHHgHIvtRtWRLHbYBh6hdOHUJJm8obq4sITjzslVRCfAiqDzJOVWL3yr1hm
YtjJyfwmHiWYRv4dNF5Jci0dBHNVTSJp1Tn2Q0eE4LbEAKzf4m1oAIHRcXHFFaFWcx1MSpNITo3i
Kkhmvfd9eLNSMD8NaKImUOHyXRkGpev5N0EzMw+O3DWpCVS+NwNqmoTreyEnGxJAiUfVDzTs03n8
EUh/4WvUw1jixCFldjjottfllLfoJ2kQ6o1nJ2oBFdGTOrijDSK9jWNU1hdBvVUF12lv6QWQzY+1
NPHqd7PH2RFhOmNQQrjL1h+ZzakjlVMsob/A2e/9hyf5H/lq+ogDOAXnuZyPdoI/AD2w6idP1fnC
1m0zj43UxveCknupFPFQE7EGLzgTQ4kaxANgl00oz3a+23akc8EwRvhqwvj2Ka1UuVLhZQeLJuSk
BdZrMNKYo2DXdboVxo1WeyCjDfY5ETiGdE+RRuBbbZ0BgXyNi352UF1f8oLBIdBid/itYFLT4ImM
q+5UFkX1iTFs+XQJYFOXQcIIF/2bvfJSvHNY6CgzcbgBqDegq5pi7Asw+ZTBmzfQdgja+qhXK14p
9FH/yW25CABjGdlWUjB11hUdcfoVbi3+fm+YkYXVS0dfygZ5iHIccP6Tjlze4zXGM1I6NhaNGctW
cJawYixuzFygGQpjATlafTCi1oB7p/QIUe3nsKHGzEtfBL54jcPZ2AMAGHBXEfjmhuLqw9I1c8nN
iB5X2RtMcFTB7tPBRZHMmXDYaF0L20UiLq+h83Kb6yFdGtbgwtvqJmaTMEpwErQj7EHK8ntkSHus
q2S88WT/NwR0lNDD0uKFYucq6ZuRRqBzC3foolpKbiSKIoYjFV8l1fCSnJ6TT3Z1WxWkHOdWCRQi
PAd1lgGP33zM984Rg/EBxCRHmf15Qisj57KTxkg5tsAwNvlJbFMG3NSsHIIzhRuCzBNeHh7gTEZ+
wTGYaNRSlc7uyV0jvejWk+brIWE0hCNzzjNRFG1nuEZM27Mj9EkwmPsyCZKIPMYWLbmlaY5Gas0f
/4Yx//QVSypGW3poF8bznRqR+XnTGUcovlX7ShsoYvzowGdEhqKSMzkcqPmQfKhwKiYS0l0pEiUc
8R06yduQBILasedN5xMSp/wDJH+nsoPOQ8lXh0aCRYAO74qSzq2MXbV9D8ELQMHLEyxOnBi+w+CY
zM22z4iO1StwAP9ytsP3hlqdy1GWmrKj4ngEAsVVgYixTTSHvadJDoeDpF3c+y2rsXLMrza0wJU2
PJTALGt+utP+r2Qdlc5vCkUNW2qHCGA8RsFZ3+JhylWI3dWqf9/Y9py3Srp5fcdWyg==
`protect end_protected
