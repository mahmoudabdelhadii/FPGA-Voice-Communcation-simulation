-- (C) 2001-2016 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
c1p0WrYTytjRuJPb2T7w1zcsFAQCo0KR9m5mRsTeeo07Uwqo+R+pAboLJ/T7VUAQCmWTIRXxDgDY
m0hLhAf9RMNk82FQM32AOtvKCcij6kg3cs+SL9dGAfNWtPM9SLzg7OkiM/n7EELhbylTXn3Vrpv9
QZ52izrDY4qcReua8YY6xKZ1sP9x9gSexxMKjNmsxXpsw/I41viJLoJRSxWaasQ8LgtgsGN3e2Ex
Gs2oNpJboaLTnKcKNq3pcUq2rWoMHLOBSsgZlWop2z9juSn4/faL5Jh6ApzhvMfZJf3b7rphZvCj
iAx5NJ9SmRbzz9ON5Co40xACsTJ4TNdcUi9cRA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 11200)
`protect data_block
FMQcjdB6IUPYutnGHRRgld7l4d8Dfvka3LtR+gayejS5Of3G52uDKBwgJ8TvM53a2eRTZyRYum6g
JFpCZSKHK+825kRwsneKOXlCINq7zF8GZ4O8czd0llLz2H+65skJweEP9VFylEzSA712wFD/YmMT
IweVdyzvau3MXiX8RmG7N+5XrVULO//XPWfzgHh2MuSt3ciZya6wUAASbJL9oGqm6u8VipTa2iTM
dDosIqmBOE1sIRJcQw4iAZGw5OPzspBUYhcOnkwtXUWohyCrJz/V07dRUmtV9x2AGXeuccz6+HoH
kb9kdLFUlkvumxvajOoUMnjcTrBQLeIFt0UdNsfBd41qTFSzWbztrYZK1iODlRXGbFfzp6jehL3k
84Y0DdI7dAhyeTAZ1U7JNh6PBQYRfn2bbt1Sm6sQyisSm3gaQjkBunSES7x1LRy4/sxShOckw2nV
6K/FwjUx3bNb1xCXAWxEg4NqQT3V7M6VGHOCv5iPSrvUZ1b0EXRPibrnVeCgNF34v9h8UCQmaZhp
zLzkd72JwcAxX704nW7WlP7hvyyujU6qYED46E4u4jF/uM21ViVivwFQWO3LAkdYGRUH+/PJqHuz
CFZ/JLEaNLDu6OtR1vcL5uHt6E8VO89i9pibmjv9MY6u5Webqp2zceJq7GtTr/7k1/rH/1fzbeX5
TIjtX0pcv+jjIxWwvLFBedvix4lPmXd/3luJZ4GThKUZy/JJt2kyon9M0F0Of0O10tcV4te7yHB1
+ZA+pqzgyjq4sWYJwoR1ClmWbCwocuBAZOqnsH7p47OccwDmhOLHn1LO5nZVtMLaVZ2SC5hgOUHG
x3+HYaVRTC4VNAt38USXiXZyKo4+pLiUAz/AQac9kPXLvP+2V48g23Ut/IRIyMlOkyVl8oqgii9Y
UyOh92ALbPlbs6dpQDYeW4jhmDUbySWQpr1BHsXUMyNdTA2GlyZ8TAH16SIxVvDb55iCbVdQ37sE
dsKEWbMrB4MBeNDYkxPxvxc3Jkwpo1iAPj1XebQ7OMydQtxiNQedGKQL7facfX/EyN02cOO2fUmA
h0kpYl801wGvB7yhTBEYeYF9MNkTowFvpO/KTkYXpTBQTmUFOK0oYiX3Lm9IHb2lrNUSmw9Xc2ee
NKeinE3fRJdqWpmCoYBtAplW7I+BPL6yTGfYto/3mRBjMxXYAF5NRLg5BKzqmA6H8CrNaTpyNFdo
z5NErtPGoh8vYIcT5OncK+lKVUiPbO8ZqQxv62UkixzMP0el9CESTb5bPh84YJfjihCwp1F9bzuy
XoNgWA9IMzWeVJ5Ib0gh6zHkf0WsfaC2G1ZPHKasn+RQF9rgakiLF3rydv0ZvujQSCJAy0Gs8ral
1yJqFgEPJUjsThbW9/oAJX5y0BNZxhUDENK/yBpCBCV4LkVbg0JYhsIzn0t0I25x1xYEXxdkVfw9
qBFWS+7ZeaVVi/JPM9SFE0OGUdpurpNaykHxv2B37Cn/XRHXEBj+Wu2Todx8MnUEjLfWO3w+zL3y
qWKdUdoUBTFbxW7oFD9kiekGy7HbOFIMRwWg0FQFgiTC0jbOWCmNF29RyUQFxxRN3s7F6Mhh/Hh1
MGkSHpOdTjtOEyO+zQejIL6hyQadDYzPfT0H+lo8xe5ilQOlzVz59YQLkjo4/KwijPxAtQTJ6JeH
sD766UCfzbsy+j8n6ige3hEZ73DQnpmCz3ZEMj39cIQBdAi6Ge520exUfvxM6ZxNoJ8dTqhqfRvD
ToqbSGMEIVDFBR3SMR4GECRKepgBFinIiDjg5HcKla/buWHi4pZpk3j/I75A4L8FfvQZz/Mv3oDW
/5hGjn41uIlZSXN8+T1he8OaiaUWXLNEWq7ppngUxdo5bkkgqA2hj0IBfUeCbOSjDMzW2HefIBlZ
og5yfNcBQJkFFKTP1ldozRSyEuVbhPMPOHWH95xz8isUKaguOdYF7FsvgxMM0uiB4+QJ/1PBo8QJ
e7FUYDjZ7aIy/AnqGfTh8Q98eRR6np7s7XiNmQDehZ7N8O5ix7aWo0MoqQ8R+qDCc9lUQsCUIB2D
OK/8mNppOefXq1zUkOb2AetHMc0nIN5eEERoXPByYPA/oQWtq9VqvkP0wAEd082SWNzVu6QVKwjf
dqR//8yQTH/wVB2IW0Gq5aoRx+P1zINmyuX47GNy4XU8ZZo0Om4uUt0mmLCYzrCkBOhilwF+pd+I
HaucJ7GEamrIRPAyT0QXTh1qoIi5SbBpYm5QRpXbVqzN45VRkZNSck2N4UOaZYPRWEjrvPllI6Ix
ofk7QTWhQJYpTQqKhiURO0M+wUsfO10RJIXQZ1D/PR6U8ryE3xD51G9QCP19zrSS/KBXGpjXvyKH
foETT7OE4Ga59TvtkJpiPTVgm0uridk0s8V3Bi+U7IvwvSa/wyZH5AsYaMULY/6c+nju6VFAX2v/
oVDKwNvkv+V/spmc/b8ZWekz+cR/zcM/iEJOzpbeI7H45J7EBM728Ogqabm/VX+fj+7kEWS1QBvo
3/YtHCLT6yL52wdYIccDjDOEHVCzEv/18ilfG4xKNJ/4mlF9Z7eA9g0zORV7tPUEbykrERRD5i11
sW80E2u+Ggnd8pU9f/aYBh+o+gKwv+4oNRwuhldNXaKrZ5LmY/PvB782CC3KZcpCWbEL25txm5G3
/6uPil7K50T3XbP+D8ft45CJqFKI77GzGgq+9ksa7nKJSobFX8+Se/N7FYi6YY8X9RuRK7JE70T1
IJgMVWGOzXhFtbALo2Pya6JypaBLQWVKG7CoPpuc3odP3tqLsJOZZ4yXFZsRPXjTsmCBGbQG4zCG
g7hUfO+A/ygveae9hX8h/Qw3uADcKgja2fsvIzPcUxrAKpMMCFmKYQlHXERw4xiRwDvEKHLDUuVJ
NZ6XozIMMopkR8/LHz7mvcxcBzBDklHn8gAUi0VY2gzhnu8A4paOG5b53std8q9bdqqhsYDH0xJA
YhBPTvt4pFedcmOX2rEl5EroU7JyXTa1iWufzcwlWl3PbniLHh1DhB3flvpQbSD+LRlou8K2gzYX
TY5KKv7hiJV/CI5GYCItcKxLq8OFwM32LWy/9N2b9PhcVjLO+Kh5MW2Yb9OhPvlP9xNZAkKNNlGY
iMt90hSBlVxQW7yRxGSc6j+hJHqtqOtCvnLSfmHUsaaaiXaV/w6o0xv9L7cnOkQy7T1fwH6amyF+
gxQey7tM2bBsaXVFfiiKr7FYzpglRy0oVLbcCEIGCedopfP45aCq1+jSsv9T9AcK99AV/xPHydPm
B/qvLl5n4j5e8+B6Y1pLAeZ70jUyS2UsnuEDEj37fNEfzSRzdSVxXULDNsvZtISnFP5zTNCOsd56
E6buUhBGpHQqDdBfU8D8uA8S1Znj3eKu2zDoIxTa6Eu1CXNN+eEFCj3BxxpYGbiTq1ApJwULyAAv
mXEPxqHzMo0slRDQSzUA+cx58KOdz4gBvYmNcu5OV6pEv0WMOrBSriBTwR0pOI9HIYV/Zroi94AZ
QZ5FczcRDfSxwEsqjKzdVctxkzyXoJ+fFw3ZdqxXg9HjgrUsK2CNB0b54aHzgs8J2E3/d4hfKdt1
xV4VfaM+H7FUSPmluh3Ra2L71UAM9zDvjd14/EpUqzmwrzr3OiFOFDh0WU3GPg8pGr2C4M8HgJkv
wNr/K9dEHZW/h0byhWSF1u9CvhinRtNIiVlUOTMUh0i04UVc2wYIPzNvZgD7473+TlnOr9+BnPXM
ztuTe1hSCcgBEFPpz82dl6pxx5LDgNMT1ODrZER+lOqw4gVXbmYYdoAV7H6rTpGTWEpjVEBvnyy7
DQt6lS/aytNSeidqPD0s4Klamx1KNu/s1QNob4t+UAryHMwPsJFDSBTmXpxWJkkghYKzQwC3pjiF
cyYQk2vE4PFZe4lRQBNoxdZrKpcSfH1yTYo3cCTa5YZowKvgyz3h5HuOlao01WxqGAf5Iwc7kWm9
aiekoYr2tJrzxh6WJgv4ma1v8h0x+ethS9q6SZ53hEbgGCaGoJ4Yvs6JriOZQr6xry2Cw2ebVvA4
OpeFaIDIva9PwiacNcZ8o3XR+m9Fyc8mkeky0sjczvwR6DxUkheMEtsV/fQ1RHmwBX2ApuPokeVR
LNEXin9V+42rU1SiP7Ydaki3a5T6EK2JsHScoIhmDkxXmxkcpDw0p3z/gp7aa4ZK/zCqCBQpUPsY
jZgMrfobwI4K51MC+GN2yA7ACFNFwpa50L/xTns1b2xYYffVW7q2/OkzxPG1YAl5DQSA5iGx4Kvg
6Y+r9w52ZnQt7Kx0mpDQART8JnKElkGAdyO1eOPUJ7HkZR9VMmdIb1+CqGN0F9JfZ38kn9A1gZyM
HVzhkyOmk6jouQAJ4gxJyHfeejQ2r74sytoha93RtF8nsi1MKdVDvaQO1RtmieC4smYLzUPwRrba
Ks4gGy1/uSQIsWf+gwjUzeTO1zu0WJqJQzhfV79Rm/Rn7cucaeOLPovU+AXFWuHfWBFJ3fdTB+0x
PTrU4NdKg5Nh21ciH8d7k1WZc3qBvXDKEIvll9hRtEW4fn1O9y09fHOquSnNVghXqLAuCmxl6rQK
J1yUVo7npDE3m4uoMWIWEGkqlYSP8weo5KeAy+QnuUlXsRyaxHVPhGgN/l3xCacmfeDlK9e0bOPJ
rbb6Epg7so9M5D+0QlA5qK3aC0h6a6D5h/w+ECfG4q8HSM+ZHKSyUlsDw6AEghWyUMceNEItCxew
AbE7VqwuS7gAj+9gIPDDSQawUJs+3yxBCBszH6d2XAmZJdBudRL+AnaMeTyDk+Vu21qXaRe/v90f
lbf5Wu40/1+cpGLYaeJ1mmTs3LWOCHtAtjWuXKcEK6zTedotVJtA+wOnrbDjrR9ktdYn1XVlbh56
1glwq9Wf3pW3BMCpAMbCdpHabRyOk71/R+ayryVZU52C/s/O2LRPWSltewH9rVRZvo/Fw8S/SROR
+GoECNK/Uk9HIk7Aiv+L7F+HXRtjuHLsB+PqkH+PY8y/qXpT0b1JuwTESWAP1l1K/nmEZXVJmNoE
yK21Tz0xcr7Yg/hzP/7tDTJwN1oEyW43IUVIQVxWqSyCOBpm9OCHduVxX3gc8H8mUokVLCpdbnrm
7foC7s0kFgFMz3Eb/zuLndsej9TZXV6mFSQ67UjQtzLtUl9lbq2CcDVtKrxjCrWUXlmpNrMDEAbY
iDSI6nisiHzYZXXor95Ds9QUEe0GBRoyVLERjV4v5+HJPyIwjZaYH/Yi2g2xOIxoK7kMhPK+V8vo
YwhgxHVD1YmKrZm2Iegz8BFaAvgE7L/P8mepDQYyV2Foo99SHcjjmnneNDe+49/PzKRvx+r88Myk
TEjd5d3lH8Wg/nTaSLarjjefi0lBfQYB7cGTH3yiHCefm5g4rm1eAPlf81FD82DO/LMbs/vzYW13
Uj5NBReZEH4cahvo4M958fOCoIPGTuBho1/Q0rz5V6H3+T+MKWs4AsA5tWFh3WH4wTDOKAkAs37k
D+BPhn44XTVEK8ywQaMiiSFkMoif1Vd8Ag/WuqmGEzh9n79EuaR1dL0oOMsbdEsmZT9u0k2Ybpeq
tcy5tt60hjG54Yp/twKzMeZGlUodPZ2CwLbpasqyDPLR02HlVzteuiSoAatS2dlYlekgi2yE4Sfw
uHNAL6lrJ+BylUWvtYagcRn5Ctv/uhIoXCqCNB8eWPy/tR4TdjEA6hgl8BU4I5yfWze7JvARzWO8
JKHeep2UV0OhN5/v+P7l8md7iR1sO+VfND9xbc2fe1Bv3pfzZ2bihHh91luFdh8S6eCY1Bkcryew
94fkvLtApHeq+aYHQezjuOY5fCWzwWwQuyNvqmR1zWUCxo4h0wDZRJp/AM2tYsIBVvK6yEYQv9nv
ekg/Du41Kk6XPX/l9XWIl+ZZFtExZ5/nyP97tcn01+kgxwhYdWQGF2CH315kHl3tQs5rYGLaujKA
tSsAzg8wvQ2dWs9U6IqRNpDOArNNDzuf7jHxXle6dKLA7PInNmeVTRL59QyWSzQxxzkIf+VoBkBq
KSs7eDABDqBvjTjWFxG+kXd8/bASp+2weKNn/IlyDRvG07ATVpNEDgDROiW/1XOukrdFUqIHxtiF
8+5aozLtTUlWMFkmDaQuC1tx6s3rVJvJku68Xe9gkby2PLAwZlh+CC/B3qfEoNbzG7tDwGsWuj9M
i4F7GVNL0TVTG56bCBaAObqoZ5GpRahITUvHutzEh9uQKtYanzVXvuqWAFEVgUPoAq5HO4deyvyd
jyJJMUiBC8iu05NYp2TCvYO+st8+qFmIhOvFNdJv2IfRFKq8aZC+3CZ6uYpc7VKU89aCcRyHJS77
AQeJECB4sT16W8vkhxqiJ5Mm6C8aSmhDIlVUV8/TDUvTOp6uhMbmENNnJgRlsCxLycL+4yTYV8ci
VHtjTtMWAGOj/mx7EMwtOlBg6RJ+S5zjTCYN2WtYIqtzifUWXLXVq8TZwuiM6CYEjnwkkutSMDrc
EaCekIRaA6aRRmufe1f2Nl2YmHWiyqyyLgOkjSQVL73Vy8sUjGBiexReu5/MCBVdHM0LsH9wjALg
RdxKjCPFFyiJi/ntqqgiQIqIYfeOQhIwfy4cqlGlEM/NMvEHEY06Ok99041NZxY9aZUby5CIbPhg
eE6kiMW+15xZ4+7Brljjm4E1X5toAPALUJxV3JaYZI7Qo1T0tjsCg8sQlgY6f3FpcS/dKy8dAJCi
e7c2LjrPhRp+B8K9cSi/8hFJUfznGvzYkDQfBBgrU2Jx4/BEGBb615HANIJcHo09QAVzzdp0TDIw
1s8A2Ii8pwOoUn30YzVEUPwrGTlZ/EJIu6umtLX+m7AH69lBTqyTKpkVSrsufrJm90lW3oIssmtv
HbpZEpFVq2jLi0bRHyXWWigvhLz/Ij00Yq3y+S3kWpLmvqnKo9Sh0xXrMaD2gIJL4Fhp7wUA/SEP
Fl1iFSJEI7XY5khUITKAVVwk5VbEUxXM2fL3CC3xO1JnFlhEYq03z2R5rZ5Ov4CWA6h7Zbj05MZd
gZdy4sJoIB5vlF8wfQt4h9H/iKlJSbsygs4MJbcFYhCqpFkgvqEaAKovbF+w0Rvo+VgHv5d+w6t7
CpmTQEkrCGTjeyMd1SzS4cRK7ES0SDqRn0ScaC0ySR9dPjcWz+Qv9qrH/9LxxnHc2UgFA2hXHrCS
Zps4fCE9ZPX7jtWlx3/wdYZUdBTSr+epUf71tMTCOLijgUhavtu15wvkajRRNZjgWEl3yoAYNVE1
nPYWSWbUMucF0dnudZzmwLv8KWCR+QIipXOz57X8PWGzGJdbuuFKfITDAXAXtzGLNlSTJVIukzqy
4uC2eILDOhxCczW1229PBJABGMrIAxyY02ZyjeUtoEqKqKU1oRdjGYiIrilt2tPXwhmiEAdUx/0C
M4LEGOkfCdjCyuFNa5lvvVOx/LLEG6ZnKnqTIoM9cMoE/565vNGa3xjCSGXy02C0e/ZzyCLmRebE
/CsN/tTvBFqzLhzKKms2aefWnewA90G4sytWZidFYINhbtRBISfzfi/7n6nvpp8P9emia3Ih5fkB
ES55bqf4O9YKCf5fX72rNZaNT11j78tp8F7ChKhH+5RKBWWOwwdZorU8Ub+bMQNFePD6Q1C+e65v
umD37y07vuvOPhdgBtubA6TJMgoRUyDafYN27613ZeR9Uo2mcafQ2HP/VkWL7fEAGVSIpJjqCxTP
OJ67H0xM1pCEkgFAOb4loJ/Pn9Er/mHI0vEMcWxMmfORphDQaeDZGVTIrbgDYZxnmMuBH90jlnm+
7/Pz0qh9ndnTwaM23dc/9ELidZ+pj0cxfsJ1X/OG/xC+224wNByiuOFBSAaFPlFXdDgzcNRVt1Cx
sSsLTuDayNqaa7RTPYuaogRBZyjfICkU7+ZSf7eBiuMCvIk8KEd4YQM8mHghpE4hfLeOFCBdbHxR
pWaI8B01hG6Bb4njXALnIEaqZJZGZjsHV5PaARInsQLlX0fc9CLJCpCM+i5SRx7rv6dov2w0LiD4
bsxwR18OBkTrwmekbJ6k9lWyb/m63OZZPxoplu2qhNOtjavSsO+zxoZiktzYbEb7/7XntjoPzBkU
Lv8NvSd5X8RtkZDLORl252dsvtdcCqbHDaVKW838oNtyMi2e7OB8kaLfRyeXfZ5LomQHLUICXoVM
3K4crOF7FMtKBucQLfn142o87C9IKGpjI2rYKcNz1AzeJYSmV8Rod5N3h4jGl+XBn8hbxkVVE19I
gix3Op655KABLLI/Hw9QYAyM6Xg/9QP/c50DuHuvCi2Zlq+uyCqnpnQ1klY1rNCeQIdsI1pK9ATd
PodigfeZoRDOcV+Zn6oOLlvmR9sCfZjb1wlazFiiC8Se6A3MY0PGgnwVjuCz13D7LsiZmi7xT5YA
bDrkhpSBfy18OpwvPCa48GttWAw+w63rmRswdCsDZzsT0hf1IFA26ihGpJDfd9ButEqqFd9bP50G
wwUPpY8uKcIb9dgGlajOr8mwIgsnKwS469YNzRSrwwoVGln6S6Ip75HI2lhHJVlYcVmCG0AWaXah
eio1k/IYgPCkklyZF20+jfp4Fo8XFKpagpN+OuApzXujwglvCMwL5wdQpnaNQ8TuUAIX9gVG9Mt3
fsVa6+mSkiwHSoKX8OxGLnhHrCLTzbXphLDpDR3BEMZCvE7OG9xcTrD3yB9YjB9Qg+Nz144VImwZ
/YoWkXJ0WwY+5CZpeI/u8kPmRvmhaOTB8R66lRo6xwzeLfc2euZnw5KzVWWmOwCUkrGm015ufxib
e9+h1CGGo0i82EhewT/3B+7e8Gj9hQXV5LrU65mxCJRSokyGhdHa0IiNStAG9vQNuDtStfz0db0h
n47NTMdk4+eM4jVkel5+LEpH9Q+rl9IDoEsj9gtq+qrxs5yMX87oifuZD1tjkxzG4KpwpsCjepQh
62FCrmteQTyQMTCLAKWFN9NvkcqsirJ4qErsQ6meDSp6wONQZ2MNGAaDDuJwwAcpNKVWEufVG1aI
Btr7Hnrs0C+uheBw1gW6dKwR/XWRUFRU0FIQ7W42CUFPABl+ixjxxabFoPWtVelz/DWHp30Kmvxj
ZgeBXGAH7poHayl/1Oi2uofohYz09TPDBVxZuOFDp6U3+iCHnDNoI5LpmJX789x9ynWIoQxou4Qa
FbG12a3UWSUDp1zZe99aaAp+8Q8H4i6m2AztdI0W/f3ZPFHwkg3gPOyusoDqviZS79XrsYzPNNtK
lOa4XoVxHcs1iG13QiLhK4jmsbjhxLmEZipZUFrN/GbSSloE7vW4rcVYGbDO+s0Feb0b4KWIAAtW
7wqERs3RqLSiYaMvvoPRMA3hhOor7rVBtBj04iEjzFMcGPnG41SRRX12slPSaDH0hzfbzrngykxQ
2IjtJUfYg4HPCW0/KVevT6G7zQ/9pWw5eMP8vtLEXKNKYW71J+65nab+uQRbG5VowLV1hKSq3Hdi
NOc036DfziG3sA1+I/MOcJ7sc5AyJOdRdM5H43TFWyYx7q1GRRDaEXnLBi2b7SEOL2vyCpDlHBsd
YWIdlwqRNiGa6fLKPdoLqRjYbjLUxN3IL+Kz7N5I5WFei7HX4yCp5bOWsWavxThfYtZDOIGWihOB
SzwxgjN6qpyzTzo0Y90d1N+d/ycDGGiMHf/CyaS0BZSVPYzjfZGjf7W6FG2h+u3F+bOcMAFRPHqf
xLLYz4GrYbnY8WKs76GTyZRdUDQjV2W9MGixU0L+vUNT3cJ02/cI/Q6hv9KgLC4sKxGOz2wJ45Yr
Rz3BbIL4hK8HJsZXGV26tiiZudjwt4b93Rm8dgy2X//7sk5wg9MOb/EX4PXspAxeyy3mcpXWwQPZ
4y0FAHh0uDr5uSJSGnefIxRIef62+M0y6z8Ms67pTYiyNhOJ2OiLD0s1EiuAmA0S4WZ1EHRh2Byn
J8qaJuQ0AhaOpCafoy4IyKQ5GUBTQq4d5DhjHz40DdzLI+Vb09hkpOeXgShJquqcqiaxcVn4fRmr
xFgillb9EPrHYfxqGh1LTfPcLfpmZRJJLvhSva34Sq10SP1OXtjHl/gUyGiCG1FS4nYgRuwSh50z
/h+ak7wDL7ph98JW5dnlDbTmpqih4rTPbPcc8d+XjDLfvdEQWwmmR0T3h6Vn3OtOkt2USHVosBJk
RQFMWdK/hMhpdZ7QvCAwBueQPSKDFfav2mGlUL67uGPSBEWyUzH6g4orJhgN0iqq5KfXGCVuyA42
OS8m45BG9Wy0pfsicBzbO4HfrkVrch83rVjuQRieezLT2C4R8yepgzQUx/xxFX1qJtnUFmU7KMLD
FuBnEUTD6h/zUgwFJkgLjnNivMyd+9rP4hmD6V/7Z/YI6Ez7aVh4s1zsk3rvhKDO6C80wKYXBvla
Ivg4gxtgLuhaJL4dSn3wp7JGku18ZRgD6mVaVeXlxoRZRnFhyXFX0ocb0Xjluab7qKLK7e/95h/B
Kbd2QVAjFPAL/KCBiHSOc+m43QRuER3UXLtjREEwh/oZRzmNFVa8+dospVGWbMchAz5gqBIKbJzB
ax3h5svYuPocF/4kIs6iFh/WQE704NH4Ktq5dCtd2drDNdHXXp0zpql/oIcTjhnowfmAC2ARWFC6
WjS0RrMByOGbSGNer/k1+bjXN/I1aFULuOJUMz8pq32C+LcqJB+PwAVCCw1FiKoaIDYRj5KSiAIl
VxDpRPALHjONmtkHJFB7pcFlr8aLrYgMB1BVz+4LY1DqKvNLNzPcNhuMyttNtOICjOdUcXKpSVx5
O9FUfAWlsy5EyzbSCN0WP/YEaX71K6FJPLof9IpNn63zYZnGUHxkYtOIZtjZTasz557F5Me7lBMk
OHpdyS5fOCjSTBQevC4yiieexLFaicxws58ecGMH3KwbFU33wSPfHYJsZFtgLrxXHw2X9k3lMfnK
ODq/ybkxcifBAUve60KCh+ZhlAakXQDDUmVr4F52vcHKuY29HBGzYyA9t+b1+om06WtXcOCpeZJq
blioapxMJU+J5JBOTdKBu74OEwZlua3KQ+at8GzLqGFCjApv11uVIYjNBR6BakyiBvmW+IDAxHmS
p6kRVyUDVU+DHO6UtjTrUeNfPyn7bSqYh+It7laRNGo/BeIP4AMMqvoJcxQGoheI3FMUbIvUO9M7
2r36Gl1Hb0P0WWAzipgDKmR7MftFGK5OWYBZ72b0HP+EhXMTl1gcQ+jABr8WDzRHlnBUvNcDWMuF
rVkZx7Eklr+TPJIRGh1MDGoCsRArO2xv3Ogi8QKc0hKxmoheSXmB0PBEsQmc+PcF8G/FNf2Ho1yn
OMg7mvy5JmpdVmvo4YWSy5WFCYyecnDpLPfOoYrRhjnOIZ3dsXO89/Osg2424HB5iVIRum9RalGC
IAkP6okjZm/byMj37GNZFWoIHkmEpfQ0QN8b+z7JmqxYYrOx9sV7d2BRJoDwoAilNIpXGNhUYTQw
0yDdOcpdiXFm2qmLoxhn6t+S/KfY94kSiiCn/q5Ol4ouNo+Orr0sjD1pf/rK+9ENeeeXpEnFJi/I
uuCcHKc+sxsNJtDRWbLsBqt0hdARGDleQz3Wh34zNPNR9bfan7ex6jaTBlcr72+7/OW5u9PgNfa7
9ang53UpZ9iD13DoVz7zMXvmf56oubT4q5r0N1jwlguSaUTjTEnAMb5FORzZeIO3WJwPsNc1LX4s
k730+fsKid3f8WVJIxT2uOOvrxRo2jmsm4WE6xspv9eu5W/OfmlnlaX5FPqkmfW60qwpJsJ8nBxk
FvPhnZ1s65HLIv7VYtoTa56eq3QXm63PrdsFYWpAIh6O6YS+4q1eEJ3SBftqgcbkk12jA+Ac5cVv
AVM1A72DqEgxFuXLE5g8BbvPl9Qqgq71Iup7DW/cv21UJDrY70zgTBeod72HDloAxJaVtfqdefM8
Uqgu0ur4rgQTpOlzIbEgsHyftqBWI1M/6bA6bDkjj9fP0JSamMTgxx66OQLg1FPy8eW0e10JfFNO
d3qZqL3ovWjGX8MTXSg3TrxYmaG2vfFKJe89n03cTAZvICUtLl+oTvSvR+edtnTT0I8PVXbCmqm3
qcVZEJyYE052QZHIdLzaxbWSdkMOTAd7OIioLiUT14Pj4QjI4CGAjTmQhohK9mZAWB4oXsHsQvMW
rBjeir6jsxWDq7n3spjVYPxDwLnB5FB1z6EZnwxRicJMrcMZgVTzYitvRhRWFvDIMQKbjASk1fE1
xQBp9kQj1uoI9uHNdp1esH+BGIAowl1HlWYkDpMaEOz/D3aDuP3aHOIn0O8n4C6I8igTlDCbJns5
mABQxsj7ja5dvOqtXAnH4dt8hGgGh3G6Pk4X/b75ZtxDUNR12yvbAPt9cnQdEcAaJXEf7e/jnxIj
NrLsgJN0YW+hQNKhEXQLMp24uT2dUvbXipWpEROtFyU3wDeMR4ST3h5O1xQmYr6ihR1IKzUDB/tp
nbMPVsXcgUUd0I5wgBuFkd8X9pLL5FmWVD8EmrNvnjc+jk1QWhmrsdafpjKrfW0EldNb8Z6aRnQN
ZpxULC6S4KocjqpIJ7QLqaFyfHFoqfxYzmqNLwZ1Nd/xE9q1lOUFM5PRHLXmiOzdk06Fhf5Dyoz1
eR69hvanCUYDgPB0reRue4btzrg32Pg9Ym7Q09Gtw/MY22zljg8/SrVLlO9INiBhPpIAjDvR/6xE
kQMCVNjp2qnECEW8v0mbQ86LCp4GAmTNwFTPY+czfqWrOINDZp8ipiG+gahhEDfQOBkHWC0lHWoe
gnRDFbufNW6U9pgfsk/9j9AJ6yCA8Mdm9dnj4Wp/MP6H40P7PjgjVLdRCSSZ4zNwfbctA+XDxrK+
RNl8uTjfahI1M6zq74w7jX6Oq/y+jYF9ZH6GcE54anzPHP74e7iR/Bg5UZX9vkbN3iBrrmwKT3po
RE/aL6v06MM6hUTiJzp5H7ja4gUyrDQl6LBmE1Ib/AvIM/YPleegD3X+nCBw5mPpcEPTZUVLlxrn
60FJ0EudizUzEbzB+8m2rrGbGNSl9ExPS4Kp4uYy3F6GD47cpcvbbCuF4MFdabPQtTInwmkz3Lc8
fYC83fjbT7GdnB0rGDejO9b2i4DxtefhO4z1hlxCYN9BgzpVymLUazcRks/Rm5jhRZQ8ZCw/2CSW
8kKnLSiL5kyhrDupKxn8biFVae8smYpLKb0ibVhw32WUTPD3W3njlscWaK+MBk08MKtKiNDQkErH
e8k2HREnBU9j2s7hVrspm0i3OLRhX3/lIB+rYYZssfUkMAlmOOE8Y96oneHu9aicSmxLTH5+QAkx
3QA8sPOXTCDefEITKLhm9iT5/G7nSUZ1RXnUd7O/S/P6yinJmSn8a7vWH6rz1Fvp+1s1pDm0cxOc
UC/9HMe/3AUE7bR+tMlVKXAAFbFfCgOcR2PKzm+jYgQwsN9zH1+jVTxJWkIBjKKgeI8vXj7YOA8Q
ryPQRDq2YXWq64hzxKIbCe5PWX1z1rCb3J4puRuL+f7EVvrDc0SezQKwiJU/m2rKapLrEekuWzuQ
zqLKmPz63M4iPEyW/x/xdyI9/fgiJJ36pRXDhEBVuvtopj2cJtiztHXJJm4EuquNfXW+5thp7rkJ
8J/BgOI+ATH/+nonM21qmvciAIr9e8diB+ZrTbaVIFul4BYUK6kOK/EO0fXNMwP3AUnNRwL63EqM
Zu8yuOexVdyfUrOzZp8xWepjcvjLoLUTaLH+bk7KjvVKPR4RfikTRGrOo2OB1NRrSJ4rGZXoc8Yq
FVlunb6VbrseaqRy5zbH9FSxB+YJO1KehLDQBtk4hfCMW4IUk/2SxyFz+OYU9ut6OjqXxPpyIzkW
FaYfxmG+RyQGv8/4Wk1+/PYFVvxAt7P/epXORcOoj5sAQgsx0FzZMjYCatcOGKwblTzrHqY6zCNJ
TGMKw8dTw93jTsfNPj4o8LyxFdOyriOvDlXUb4ALW9tMvj9jRm2ubTB4n1sH2WBwsThaRfbafwWx
6siIIklT+unEY/yx22zCZoyDTmzakZD0kkjt8jG3sPVgfnrCoyxZSew+HUmu20fAwd2bzkaPraxt
pdJ2vmvRmA/o0qqdK2GSNyVAVKu/RIbk3rGIlGK4ocf+hQ4LkhbT3JNb2yrXUxRuiGEjW4uQtFmB
2UMQ2L48B8FSTvMnqwUJLueETBNzXPs1nQyV6VP5/YS8QmHeV9MGKfeBY4znn+P7IMF990tkQlXQ
kL/ewQ+YH7cUpPnrF35csoQjf1vQafC54v2Q33cxYDgo8jXBdkqG5j/i2QdEuLES9Zt8kRSKumOA
47d3qLg3DtV6qOCPR5fgU3vceYSpz0LHu+r2PmX3fj+DTUWiY8cscJeYVuRomlESEnpGkSulfkJs
shx0jX34SrTc9v0krlW8Ziq7XKpKxhK4H3f16cYN+EmzCKBRp21X4fOo7nB6MMeCiqJoXK2HXblP
5BVFJnlZ/LuzxlMbF0vkaJ5CHur3oMO6wocv+3gnQ/eGypqQuR4A32PVZTBv0ZUQeC6HwsKUveG6
xTVZqjW2bYbR+UoZg2zUL23MOivuVNPL+FFthXGvdvjpWZeN5eHDN/4YvzWNfg25hOJBfMSbf5g4
wr/t9c4/4mtJo39jo7UrkszVgQ5oBIBrId5Bz5gKUe6WDAC/zeLEj0rVVDbl32J0Zo7RslNXDMk/
8L4DighaKKNbqQLbz+9aHpvx5Bb6Nr5sCGbpRsxzoEamYDZafaMUWu+JDExY751oSf+gUTX1ughj
O0J14Pn/CubZh46l/lcnqd4Kqtt0xPJ6sT1b3poMp6UR7KP8TtbTdyCo05ZKjc5qjolQQiLtf884
N0rEOHpPVHfoLLzXa8F3wUUXrCk7CiwewAeUZsmXuomH7E526VyDabZN92pAGiN5jRk7n0oW9W4C
HjJQLvsE2qrBYGj2kWRuVbjhSGEiuDgpW8L1nrIODFGL7JlI/Ddn3YH1W/Q0WMrdQ0OQgHhIMZJ6
m7EmsJgl7AKIQy8ojhsqIQYeyqudhqN8+lFxDw==
`protect end_protected
