-- (C) 2001-2016 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
syCG5KXvqUjLBtOvquxiVgpCYF2oO4Ep87KGcpqOa/oB1/3ShRh5trzaHRktbEZht+xFUWDwM+P1
m2fSrVkm8pklT89ZOkW0Lr2gOfMsUboKUBC7L8jYeA59kpr/TlgQhn370E+JxKeFRPWjaiF+c32m
8CDex1XjH0N6XNly0Yn8O9wkpFDn+FwbObTPWPRkOO1MWuejClczuImx1bLxAND5d8S3C2NmbQ2c
YxhxmePFMpvPlLfF94fXoD4IPHBr+8La7fz1zlKngEKXhnXnEG7l4GtUqub3tBpAv5fb9T7rPia0
9dRaMGqwqoBMr3XKBhV/o7dI/RSBSoSxc3igMw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 7520)
`protect data_block
7VBXDV8dMB5eqWXdwVmEhBb09+zJGha+cCXguPqqJ9lOXfbkA4bFElTOun7xa3WcrfB1gYLhWJvB
XpjsInLiyszulBBiBJS/MOmG+GAkTzurTmadzl6CwVrS57Pf1PreB7QxpONBRpWQasnlk1OaydWy
VD4UzjyfqKnKGKP1eHlOuDjxHH2hAv5BfQl5+TFADhsaPLK61AwmjQD3sqgoInfMPQsBwcI3zJBy
EOlL23NeqlBqChDLbmW3UQ3M5NDFBdT86livlEQ37tixMBxePM009WfgAc2stV7UsfIShq8ByKlY
nse7yVHVMwa0tVbiYNggPjLkWX2xEMDmK/S4dAk6tbCiOQj4AQL9EPewRt5d0GRVu6B1zOCH1vYP
pc0jrLiQrmYvsk0QbfuSLRgRCZcX3+Zt0AecvaAIT7ey96Pf5XmphZcNYFSLBfyrVXBWKpm3A4BV
28U8Er5V/JpwuR6DIfdgkF4u/5chy9pcS2o3eIXtBZoUjyi+rCbw77zsDQMHA6FHvzcJd5yYsKZN
uMLirKtIjckjWfm/R1io1RLHkgGwDTu4sKDZ3sYrBJAyMyjr2cE44Eb5dAH+s0tCbealSa+u+jL/
pHpbhl94lr6Uyoe6Lda8PJNjP0s3Q+Hh9CIYi3YRs84mXiRKT7sMSxbjZ8UwzE5A6FMq3mzrO6Xc
/OovlwhAFerkvGgDnusovcRf+8VvVLJUexZS7Q8I+yVcif3qRx57KuFh/Wd6pr9ky0N92itt6xnB
uyOEfH4l1AsmsvOHU7Z0eexZIruvhZQH2jrlP5O9nYMweNw2fcqKwy6MNrBPBu5i+lR6am4SopWb
/OhYvwa0V09q/Q6EmhiZoTLYJOi1uOsopSbb0RqMTh+0KUxNBmSL6GKX35/vgjjABMCjTSDLZMG3
xnPc4Jaz2ZchrYuxRkDjJ9cg1gjSOaSnImryETVK8TGAydp62aK4v9rcsDEYxs5CMPV9yf6lpZYa
NG19jcmt12ZVuS2/tRoOPVk4vTNRahfzHzcKJQdBjwE8TGbs5I2fGCfPuga1Bzau0+vUhsyygIMn
fVVv0yuD1dDJs/9JvWKTdOdYVpPNZU18rtTDQozCx0NMwvZoMfhzVquDZrPWqH12WW7cApA31kPV
ihZW729lVhFcQ/K0tlvktYQBB0dT5cMB5CUAxuxbNmEZ3FF4zWYaxd5N4MDV/5jX1J58nsZ13xyM
gxYDCJ0HgfOMUjsoEltuDQX4wIZbJpIPRy4xGw1oS13VL1AjhGyoE1oQCQhrSmPhIM4F8OLEfNrr
miGrW/LrIHOeR33i5/uUPg/Yrcpi8Q6p/qK1Nh2IAyj8idyhmyhNrQXtLoSfMxGsnV16ZJR+iuc5
qVrnon7ErhM+060dB8NSIaW19sKkBskDnU7G7nk/XLcE8OS9RJJSSl9tHYwloXlKfKpAH54BN4DZ
wrKTsu7yjBUgI82S/CgUO1PSKNqmn9YwQ6ox6y0c5Z10D8JeTgTzJE03UonlgeUMdLRsJBDN/lKC
b7Kbbwg7ZkM+mEdKYgTVtf3+CNk62BSqTOEWNVQ8A4bebXqMgAU73IU4S9rXWVGzdhoGbojm/7ze
/C+L2rwRheT9ynKtslyzpUxdr52LQP8BSM1pdsIUw6EwAu6oFS8BrMnKN/XfvbeGxAEERnXzpBJU
XZWcfHZbmeGfB3b+aaREZfqL9SCyC6Y/wzDvYjY2fDKE0EVKudJMsuasVRnsTw/KkNMAJkOkkPQr
GAC4S0rTOICRsLwsith9K2qsNCEwujwqFUZuZ4uL2J4K4AdIj/mIFbRQONjVJ5+g3z1OpKR5sMKv
DEdy2YvcIvNRIwCJThmD1pZs05pdvf6srYcL1csLNBeC+RRo4BceUeIfBuLmhauZ2dB++xz2jsEN
S8Izn9qcut1fJ03L9F8wdRntI953gB0aBv4itJBhLN4CrLfR6e0BmMFybfj2A47Gb9Q5oiPTM6D+
ajADK2geaUKkNG7yT89kC60OkZxaYhrSU5BmOs0AqYaBIBf+pkyq5kr6/UZuYq5S0WNanqGqV3dp
oLAvEgLNxRLG0381SrTpowBwpaOwmTrPpBj5ZC9neatvwlovbeuyl/rj9cH+iHiYQZVKC8BQ0fi4
ez7lxtXJvQwyVdFS/2/45Fyz0dt/KkUv2ner8PFpjTM1xRMEhRrpWbzE+lYLlbWJZBdtD7WKoMP+
g7qwoy429wyR7d8X99ih5B5Uioop4RKPSspRzaalUanrCR8QrDE60KNCwHZrLHIYMhUHirH7nQ1p
p493tSbiBg9Vmg1froP60AdzzkIijpInMbleuP+ra6U7lGKaHG0fQXKgCGU4uyS0+v1EKm/FekrQ
PRo4/K665HPaQsJmjktI3/tUHrgiGcOA5n2vFnItJwXXeQlUpxr0PdGmRlH4Bow7Rs/6aYXT+CAj
iCoZBkOIUlYzzqM0V6T4W3KQbjQojgv6qIarwU/3sUcEhntSfl3LfVHhKkou2ZjbQEbt/F8jjf7L
CMwYzIrQD3UFNKJcR4wUc78k3bmvNzpTqQjENEDk+ZDn7mN9yieDD31S0cm4C2zzgikoiKWhFc0F
ye3LH7p4qhZAyGUSFnuIK0Dj5BJgNFWKUit1W+o6XrdI+/+j7y1kjankkm1YNDyw10Y4l5r7bUh2
yhsIKOZ+s0cuTfRj1tT0CDy5YA9m/JUSbQnJfrMd7X2go7ZZWKTmvL9k/uNK6SxtHWm/2dzF3G2c
mzjgkPgi+o2TBPI+xQMd4xcS++mMWOmJUStEWYOXnKaXIHZXU0JN4tPfqk93iiOlH+tI8LN9p7cg
gurr86hilxaMX7yYnIZcB5d5NJEj4IUw0j03nzGKHEdu9JAjLqQ0C85Rv95t7UfhDG2yVSCVZQeO
zRMw62WbkYCnjO7h6wUS10INmB5bXlMz9GY8id5rTqwt3NNV+wihJ1nxthMuNFW8JOU3wbHZoWH4
i20dEknJE1vWJdmm3OunASVGCWanFF23NtJFi+icG+r0hVuC6kA1HDZ7ooUEpkbzVLg5AD7lcKP1
kh/55G4Y3mAUBHiYBe+gUczYYOig7GCopRCZjWhfSZk3+j2Lcad+sqZavy3/1LTfYKf3hBE0jTuY
iGyXJg8Nmujvx8wBjMXZkdYM5TOxcd0IeT4XujhA2teZRF2E9tWyGOJ/6ysWbAUMz9+vrH3IdQiE
rChE3dz8amAzcdOOpRsHk+tNfkLf8SXpAQOA764qTFUd2xXjlsCZoHoqHQjqk6zs5ZguO5NI+Mv/
j1TH8jkDeh2JqMcL9SZ7tb+pwIo3x9Oby9Kg7spNgVvkJ+o+z/UDR07a/mqEb/1UUT9wFmSjbMXZ
h+eW4qkTw0XAaY057qyEI/nslzAZbB8Oa25uhPuhIIIzbWgDFkWTyOjMPpZCQHfoEv+0CWAl2hqu
Vo5dd7sOZlmxnZyqaTEv6ZFGYlFFiXZUtFWYTY0L4o07HvvLUq3ZuODq6QHxxBifeoMr5aooD+X4
jFYcTFaefDjgyN6FEwIloEKUKWg+OcE8e3usgS/QB3LKMEtJFnrK4E5aEtF0mCBlV+JVmkCkvLov
A7E6URdrSQI4N5292s/aomXHVhx6pJF52GLX/iIimR605pvPgRS0gCMq76Ziwr04oJVVSsVMrwbp
BYNiI58sfoVFnolgRDsURpIgOCqyJ3SgWmjqEd/mwXzBDVC2MKLIOYGXq7VJKtt3TJ8k6+NqSZS9
R7Z0Q5Z5YVyD+Jf3TZjmRMkxrom6wJJMPRxddLQ4WzzusDS2gWvqLQnk7m7pI4XemyXBATtwhpnf
g3nGlTFfmpzBqcLB9VaJ3x0mKTOPb4VtDQCDuf+3B9Ntr0zg75GqXCwrAcIAJBeirhy7VXH9GrCK
tTg8WbmD6g8g71fOyl9U3g0iHwtPumLQbxblTvXhtVoX8IMT0GJt7pECPIrYRHHmB+5XNOsimTp3
RPtJLoP2THs8eBMh9sUYSoVYeIOfMyRBOQDun60L3dkrENZPRDZEJf12ZolXFsOL0l0Pd+Zv5aED
z6sgPxZZE5BcaTHnORlsmZJjp/fAn5LnMMLdeWSzrkoFDM77yM8xQIru4cjCJd+XpkaKK1x6sbu3
FSRLe0LWHjpmSxRZCCShZ7jZ2RzLwPmTgTDmsZ8a2YBwTYJGcyswQQeMHQ9HMZEdfOey6a02K9pO
5yZBPzeBdnwx0GlndDdkPChazeTtHcvdIAovXPLpO6GEM8FMRmehAHokAw9EvVc4s0O4t+aKUY2o
dmkWIr7GzclJOum/DzlMTqqrxFK2NfWVpOc6sMZslXJFwoc2q77Hi1wltbuLLd2ZPcpmL7O+k4kN
IZ7dcPfxe0btwNRkW1Ja3F0fyKXsNxRNCiOTmN00rcdtb5tvqdZpdzC7G6lzqOYspMJUa67aupQD
l3/7k2Ugp/dy9qVUVAMTy5NHZtw53cV5IMlVZlUBoHyqPZqb/i/9eCSuQF1mFeSqJVLHluK1kqA8
PwMLcrs9y8qhYi4QzNosI+JQG0f1KipwFp+iY9q0KMvyB+An2LFiIKLEnwNcgyDFSRETm6j7hKet
VdXaE8VjuDiibsffWqhvmwTACC1T80J5rAbsFSqTZYDFMoZ0TwtXBAeU7lMKFoH0S/txzhkJgozj
0otwmh97vCRXYZuJiI8LUPq4S80Lg+cNswgXefK5+Vhfi/s1hHLirEiVD/ulCd5Fsw28aWvGNHo+
xRBNM3Zup+zwnq5WK1TaO8DBaUW08poMpRoUM9KQucX+RMHmlpmX13EmY8+LWuWqhy9i3O+ahnn5
7fWD/cBrF0HUbTKUEnn0NM14e9IJu3EiOVRrsar3qTZ2v7CU+Z+aJhRUcdDi4Od8UkfV8OFGh6Zd
A/U6aGKmdQTIIEmmSctskNDJyyhiO9WCarQUTgZxJYVS2WoYoPTFbbUIgSXXKBOM0eDBnFXUc70C
TYh89ZxwaBVRcbY0YEON6lv7szx8WOyBIxImL8IvOPPLQlfKfLKnIQ4rl8ak0CRCO8KRbx3ZJiMe
AYvlXlafsgC0zmcbRplFnS/HhiUE5i4k1shN+qcms36OutQY5aMJRhh54XRmdYbD7OOPJsTdqrrK
K4uHEzAdU9TA/F3c8XXp/ZI+Qezu/ZIbcOvpL1FFtc+BvBvsG4EUwxejoEIHUkcSQ0fUr3krFynQ
zVz/kcsKI0gbaqCQPQePIMjz/LLzv1H3hQyJODSfm5lyWTbP3Ois6CmCJVnwTkbn0VG54OyEu3CS
mnvVDGEMXwL2L3BIlfPPtvRzI3BgG4F77vGpk4z6xAYvcqwOW+5SrmYB5l/VGl5+0X/0C3BYIQmj
KwBfs4UpQdWZZqo9xxyjxGZK4nQ3GLFIU4wVcOjHyarXDyqZXGWORlyYIKdaBOHP+3VkLXFNrY19
bP1uIlKkXwOYmKlxECW+h++fSeJ0mqugyM2sH2AYzef3wlI/UD7mZW/fwCibEHevjzt6WycOtUnu
Lgv6BEYg2RHsnSkaqL/vv1NpcyZFxVA9ed3sDfAC5GUG7OqWB6LDHPdwEYfICYbgV9uWKot+zIBF
HGsqCPdUei4TtHvgtOvJ0i5SaD7xOD7IW8fNSv++4e2+g48DNWuYLPXXBeaw1FYkUg0HHOUVzsFj
LKNFzCk2jZrmVgWxX8T1z7tVD7/1+oyHjlJnmyoEfOQpJVLe63JeebrHimBO7DKozPFEp6UiN4dZ
jMlwWWOuyVw8kWcjwAZ+VK97zjH+CtKbSpBSef0JjM1ZwH1REWPzx+b6oForC2YqnH1Suj7qMir8
/7ideIZ7pHuH9Y0izDR1Pt+nZXbWmL/makyxPg005LZ754LuzdOLEIG1yHEsyQlnmBeLc3+Q21rj
6gHqnmnziHsPMwSxECjTfCcMHioc0lRo2NIawyLD4h1bEC78AHvIUatI6tAy/6FxyRywckQQbzH4
Vg+4113RuEhCgQdQiyhdXl9AB5DMt6j+i5dMi37qPCirX1/Wnj/ZYI6maHPoyrpMbN/DTqZg5+fV
+QAYSwi/hRw/E0S6+Z98knSa4J9+jLEpdvxtOLn7RdsEZ70Sy4KynRqa+TpYil6wuMqL7l+5SKW5
jQlbC9ny5z3oHbuzMu1Oa/4oBpzUaH3BHKGDX7Y8RZm8ednhLufQB+3m5VaIHvOxZVKTPf3eLYgW
KnwaQXuxqKEaUv8dKU7cWzuDvbbN/u+aRClxlvxKrFXfy9tfPzvHPh3EaMSl8KRhCFUr4cWqvhN6
sT8FpriYc2JDNSWFfYawitSg4TjzhorjvXQkuoP3CtTvmGjOvy+OMsshiOlMUuHm1Gzw9mt/8akK
eWz8vgfStHviycMy4FbhBU1ivfIqcDRFjSHoLftn8IqR1AX0YcGIXzorpeBsx5fU7A3RWg32ecUP
724z7/0+Wiu212nA0CDk6qdWO/9nU1UsveOli9QuGysYpmGUZo5mlT/FTflLsEUrLURirt5Mo7Xa
4U9It8uvvkFQdPAqXaZHjvbrmXr/VSz8cCndSJ11i5l6jQzz4iiP9XvhKWhJLpuQG6djjUy1lJux
XhIfzVl/aaq84kwJ04HKMqo/PUKTeqbYKGZMeqvtAJBfp9rBdM0HYlfbqqJI1JK5pMeE79Ol2Ql0
XrUSuwLDVcV1ZEnEdWzykOeA+J1lY29Dn164yNQxNmCfjGAKLfoKNYV46xYElQe0StpPfR89EQ/w
58VSjcOI0XvpvKHMf2/zvmQKYprXJ1OqR3XwL7waBMrV/kQFPETRi1HjUCfnAtAOlhuOwJ9/zm96
fCAAQSXerjJ3BTZj5QwTu5V+H+73NistCaf6ovcvlKq3lKgGj5P0ELXSY3livcF1hdGsl3wdlfSA
5jBL8l54b/K238LtBjGhzM+yhcH8Ahx+02XLAsh9TpHeN20eWKQu34/zoj7rahhfaDllKChCqx6B
zqQLbCrdaUbDdgdLYxGTb6ZSc6EmHK0McmvfcktlDu+rM+R9hYdlBBS5lBVzBfzef+TZuVqWxCtZ
Jo2WA8MXUJBcitsnipjlf7pT3bpfDVl3nw593OVii89RYeA2KrStmtfu6RrKVB6hvvVGOfPvQQPg
iELfwqKGKkEmaekU+EsWZVFstnNmZ+h1VzbIGonsJfvOHxhueYjzInLHxjHkGW8+CZ5M0kotVrIE
JGw+vXtCo+A7QpW1ixAHjXNcrlAej8syKwLLfMhKjjjO0w14DWoyuaVO9RBDMuiRFT5RNS7cZFG2
YCnG5P0/gwoG2PE9Js/PlZ6uRHkUkXEbwv4A1xA833LP+V77IVfQn0ne1PjrKVlIKRNqarHTwYcs
QB7NLpLEpJ1hr1CAW+lEqtYqmW3YuVAJBN8BEB1HOPgfS0fPN2Ef9A88ERcyLvjGjyKhqWADuwkJ
+Huxu9XuvF9nJQcnhtjndbbd+WVbPoQlpbrR62iCsTFv2rUHspGVK6fcRk4KQvjj1sYgXO9+72hI
lPdWGIwkiZ5FirYdwiDEcCrfflYknRfJqjmzy3k/F98OPNZ8RQx/ZOsgdNpyi47GudhYfeqEVF2J
X943VGha9v0ySLAi7VSwdtNGrG6GCuOOqO03CVd2H5ZowQL7XsFVdOdqFioYvJq92N905f4yiu/Q
viju4FyTgQvp7IeFBGYb2mW7Gf/1KQb5ndNw4qxYQw3/G5gg2tyd8A6TDMcsatT3yj8ZEYeSATS8
QEa2hdSRV6hTVFJyX1gxH4ZLOZVgRXtaP94Mj9CihjKM/QTgNpMVgVdkkkEKsN3f3RJX8OrCcn+m
XVeJu3FLmSZG+Wt2msy+S7KjwUdER0uq02uvynDP+/jLk2gBDqtOOJx5fweF5DzlNBEo/JhbA+RT
8WQQjy350mgzgZ+vMXqQnIIXbIovrtYhD60klnqkIoZPI6JXSm2FEnU0iZgQW1pFmemY8R+NE9nC
AQofEdGumj3yr0AWBvDV0z+XF81QDOlOfjuLxt4KBG4uzZ/nqBmNYhlAHu3myNZ+XEixIGC+vh6h
CrhczRXB9h4qnTu/CcXYIVr+pT+PDlXkISCNyNPv0Oxf2GlTbdmVHOBCP5/fw98FpXhH5BKm0eCk
xFf3LwpXEqbBfUOcvdW+POnUPPXMJpwIrsBnOVBtZGEy8ZtS8sjzQ6MyVzfwCq6w72mnOO5GJP1Q
JgCeHGDkyyHo6UuQBOxIZZ1/VGMhZ/YyONr05f5j1AHctcjRDUWqaUILc1M7I+qDT6lkv+b9YSza
J4PimzFuPmAipB+OBP2wyjBezmNAWlkq5dNUcqHBziBtt7eXNUd66kVyw9oK3R7EZBX8+mUdNJCk
Q4Gmo4IbQCJ4OFcVgYlNx7Q7y7HF670L+dyx4HcqAHUoKbQ7wrj7nrH0+yf+kxkY9gReFXcDur3/
ot+NyvXbn7jIihcipSAQerP4aQIFKCDxT2n9dg9qQ7iL1qdeDGvPwpPdqG4kJ2Zp2/57Ndy4RRD0
6Vs+EnHxq9TF6NUA7cKu7e8GGMqDvQF+b1EhYX8lFCHIk6pdMFX+ZGHocZrowhuMhjotFhgWYUy8
1FFRn7qvACgjf5mi7WQkkskyTZNQYmj2b5lzIFvTtv+5ADemh7RgytmCxNLKgZa4D8Ut1yUKJrE+
fYxfuGpYIPFWQX6y3Vlgj/NzaM38PF/xmSfYSWGFws7FVeQhXdYFQI7YeddaZzP/471+LZuCznDn
CWyBtKGQZ5Dzi2Rr0xCd6811AoljXfrh4G3m9eO2ScQQwhurdKugTTEyvKEHT6ihTCpJ35zlUnqn
OUnPowdDFEzKJ3S8Uzm+yc8LNYKlLRvD2r+TRfPEDc9mGM9cgkbcIhAToeSSp0YW9rl7pNp6N7Eg
Zt2twJv68kJviDiMo6Qx5OpDQVeyfZyadbM3SW/A2uJd7KcY5SxpFiaJXAZaPZWvqRUG+Vf2+a1H
tk4erOgo8umhDu4Af6GZXo0iK9VNvKG+YwsJU9JZfcNkjewjy3/cwvRnUzLC/1bWM5t7Jgk99qgc
T5PIi3gDjzkk92Bkzlb1ZKq44IbUjT8Py3O96JMceuaKMK1w2YT86cs/BI7kURvCnE3VWx3QDvvy
tHy7Ux+3TNckpt5dz0dyQ14+3yA2rXqqLEpjN+x2UdvJKUQM8ogEFWu9YKDJihfowo+YYLW/1WfI
dCymjMUdg7fZ+Uul1aBi04aN2U3q4Az0T0UzFs3iL7XolnhPeO34OZyxsTk50WVrsfrp0GAvyJJu
EsyLl1rE/IJbWkG1u4hIIEAuWg0u1OBmRGVVmwbJQW1On+aiV5FiJGJ0VEbZPDGskRL5kjtJ5/jy
toI7XvTxPiEd0B/3t/dF0hqfW+7LqI1RLaHtCu6d/6eRMfuvVqagCBYCIQftbCBEPbSAbNDIwebL
YyMlt/gB1+xqyYopQ5qRbwg2aLn36ZV9BGkytGfVgO0qRFQSE4e1+ly/NOWGtw540KPhiwVcVJ3A
9ycj75KpoiTtm73Jd0/sD7oUxXnelCrWTYWRpbfPFab1Pex4lPCr6FPy1eyeA+pfEqXNeTsVlm/3
Fih/JUw60PgQlb+ikTewdfGM1hpJREg4+MhHwqt6+U6pwUwJwILQjAIflEmZli+9FI2vhMiQmjMg
UFo999ttOYshuk9rZXB2VLE7c3V0sn6/zawQemaT5PjQ/Kzivc3YPTboEOZo1NbVvJj1CvDvl3u/
3Z4sGkZpFapY+zrMIeFEqyEbDoZMyABuEiLU8gpZmQUvPUmqfM4AZtkkPEDh96fiy4HmepzW4k2k
+aGGWFMf4BOdIkcscW9MxvtyXHgvxz4nXP5OwieyePkrhAyHj1DbB7khskEt2JY5odpnwL9jGlQW
Zf5F7XNxxg6diDegF7lY0rNJ43vtwmCOthLWM8Kr0/7jgfgoCw8Sfb51JHBEQo90DbCoyOEW3qY6
RllRk5wpJ6LWskl37NG9B09Q0yZOY5J3OvzzvoA+5ya6zVC/4soXX8lCQrIdnP94EcJyv7C/57Bz
pj0d6B+Ii4CF00s/gtYTfF5G40+PoaavFqHIvdPFz8emYIxJRlSdLumNw6NIL1Nx0LB5BYA=
`protect end_protected
