// (C) 2001-2016 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
eGUxokMgYb44G3w2YS3LVBoa3eE8+UPoZkIPVEVbo4iailf84inAi34g4W5i3FDCCHX8dhg//qqr
sbKT3hRxnpGr3zgweDDoiPUJa+7PUvigYeAnxgYhKqCb3joL2AND/KODz1wF24+UCzc3IHN5xODS
d8FuwMBt/UxAy0knTQlL8fqCoJtFn5cEtJVgJGngkQnisL5bmvuYK+gQnjw6JprKoburK2D16F1v
0CINHfSaHxZ3sfW41tgsvR0w0T4ElfjkbH/F9mD+sFgknrCp4aEYbq13gpXN5yxPzVaP9UQn5bE1
1O5LYZ1FlIgDHr7rmL2SFZXpbe/brWifdkeFlg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 25040)
S5qr7Mm7nt4mJNKX74ATkjayIBTfpVLG5o/cxKvowUVKrQU+iGA/sRKWaQQhu12xLwFz2wMCjiRk
38EYKombGmorHOJRiwW3q4mI7gilio5YdEyna+whJbBfmhfVmnvNuO4sTjNbwhOrOpkOjxFs1Dzs
gARcr0oY46/DP3/HEV+Fhmywxa0cqctjOW6kleE74KbpgWesPmIPo9f2GA6xCYBDcihhq4rMTvmH
o5btn/giA32TafJ0RywhurMws0sM1TBGDdGai+A52inof2w06iL5Vbvwk3ea5TT2Tr5qQBT0C4ud
Hy2zILmLBva1yfuxg5LUtBMHIwAEduyGhzbVChaELDcBzl4V6Vv328KAtSGDNSxP3i/Z0Iu8YtRg
5dyvYqcspTNzeeFMP6Rm4l54SPrwBUsxG95vvIcwcZJ5r2LL6xQKMNeUbyrlU/Yiua1RgIRR9P2R
1CZcID7r366fhg63LR+v2c3WROBA/vAWloqIAPEbOqXglL3HDNsx2nC6qtvPjswWtK/950bjcOlT
jFFjJOr8oBRAX45ez2RNNepTNLl7Y0bICmWb9LGCesshd7BBvQ5Gdficc/pxPp69CABw5Piv1FMB
ihnKE+56BA5iDWD8T6+yzBJ5wkvYQmPJ0QlTFEIv8DHQ0zvQlL3ajQaPrb0D+yQQbZPHn2S0b1Dt
sgP4NAa0lgZlWAhlgRrK3GCeZgF6ZOjYhZkMUlcr0tcFRQf4GZPN9rlivSeBuTPJqA5yBbcszYE4
iyB5l9cWubyIQpnib2MlEIS6ZYGqNpywJL6SGFwe2fzdfHEcdglid64BBTosJbRDwOfE1qCNfeRY
nMzJMavUq4RNCoh2cqGCLf7DIJedlsDjh2JTgv1kjwmaTzhhYw9YZyCI23yb9G1ICsvcVOAFPKkY
y1p7gDajoRKUohztvL9jD0UrQuHl74a/BZXSPthOmnsnSx0ktHNy5182QcAjGKjRfz52BxdJNUf7
EP8Gk5JazK12BwBGz017XWJ2WE7j9JGDMitSsNRgZ/tyMT4xgP/v/EwtjUaA1PPEVY5AxYASpOD1
n2gSG+B2OCRiGtyIgASLoCl1DxyyWmV8xX7JPudKgHoYJLV7q75gb+uWjAEfRRfVVnphRgwfVzNG
rVM67gVJeCVy+VrtvolL38wHi+PpV+Qrb1XMLC/rbZmkbCPjElGOkKD1lFST2S9i5J/6AZIyK5fE
n47n9AdvSuwhB0HHHIt+4UfLNsiGghmJoZoqyooE7yUKoIYtdwe0Ys5pCl4Bfl+b1yzx4jO2czxc
ODqYIPdzbKi7H7ZndnP+GVo32dA9tTVvk+ntNov7ftOnDVCoMlS7sjh4ooXlMsUGiZWICbRyEIaz
E+YcokOljnum2krWrdPXVxLupjM2utEK+ekhR49yn0gurSTj2E9uUH+D+txIk9e83WD09A3GR5k6
+LXxJLSKVnodeytiVUneMPMCXnvExE9giS7WgZ520Gm8d2lBK5bbezSe6aVuz0GCDiyaaZOxN5JK
qA4Ww7ra1e1j4af55n8qtna3zIZ/dyEP4K4J5pp3+aTsHXEF000wroc0HZg6JEU34o0KxGywNnIo
RTCaM9tCf8XyrLL2Imv1YUFb9f0Uy8oaTP63HOvbpEssTJZFtqbdYnuPIqRP+4Z5d2bLMMW/IMAv
hPvuPlo6LjK+ccnwB25nsbcoxNMxGzs0sQvTP0hW/MWb9f3/z8E1MBfDumj2MX8xWSBb12AXCPU5
e7qyKGUaQ1RcuNuur8d6MNT12rrth8NbTyUOpQ/RPfCsI0C1z60nEIXJhk0OGy0+Z4/oqVpWtYpK
YlSJhMoDjWn4fOC9L+/T9VS5ErOlzZ8/mClnEaZ+Z1fNadtRorbC1ELgRaAMUOCBAV7kenv1deew
5KjidD1zAh9KNQBjFLPBwzslr8IXbrfgT4pLePEo7MQICRspv7y0wwRTjMvhpvOoVZ+lIIWLfbef
8gKrKBpBj2fK6QbFk9fVWUrinkTZYL+SGg33LeR/MIqigNSb0s4sIpPds23RFipK1o5rd8lmj3hf
XiMQItFYiapAg44eSXYVKXxSJPvqtt3CDF8n6su2ppf6qtUurliGATUUmwj0VBKu4ybE2D9O/+MW
wrqG9RbzIbFGbKt+4bsibh9pvnIP4fkITPQcbhoQROEQltrff+eEokqpQOFf5VJRT4mlB8QNWSCn
Ps4IDmCsoBkuKhxxUi/Av/0v+H/ic2Ht1yAG3FJfdUeMKhKLXZgwk2eVJHwuREwdeIn6SpMZnOk5
2wl6EWv2CMxmIC0wN9k1zhOnNqlTvKFm7eo65+1zQtO5AxfLMKOZS6wL7MY6RdP3jVQtKQwnWkul
ReLXkYqd3uoQNZBNFTZutk8a75Fv3BR0QvENkaPvFcdQCOpM9yKrLuP55f9K2alidxq9+Pl7WpJ9
+WeafBTcv4W3JxVePdN4eGrzQxeFSQrUn4AWlljkyeJyi/S+Nnm+W3g7dc5+Xv3z/aZ29FIRtwdG
youXcVOXbaCGLsVKJ15NkE69YZZLhcJDdgVKaemR2eGaZTILzzEZoytPtwseNAj8B4j8Wb6t10G5
OV9UoShJtei/oRNpJJrsk1fnonGrqyhfDYN/SnQN4VX8mkalHcgh9+zU/IxrDNRBxWLpW1lJZWBD
0xLyouY0B2LEanjqfhHLFZvGX/BY0+GosTXsry8CNMT7tKrRkPtWXnvP1VvG6yQYoTdY/GXPOIeT
0oC791TX88x3ZMYvYlQhNDqnyRkJgPbHCZ9oPPzQzNuicDzfFohakYF+bXV2ZjkNMDJm5fAP9Qnq
ZYXC8AotviEQEI5uFKCZ47T9V14Z2HYGbqthf3WQv/gdPxnPgXV6DdKHG+BW1bD0ufxQgipkoPz8
4ebS42N3b/N3NvScXHI4M9ZZtzlhQo39+aDv7nb0yZuf+v+9nXMt91ihQjgc6X7PGCfRWvkszZUH
PEhdaAzX9HijvrUKjMf2ov5o/EDJVNyoORXwxExJ7MX3z2w5zuOyQ5VloSg+EmY6WSwUOgm/UMVd
Jfe0taCCu84sNvfcLg16HPi3Mr6EQ+Cq2C3Tpd3kBb9LHfxw0kEiASHO+0O+hoTEgC1wQRnMb9h6
rejHY5LoeR8a4SKfmj+jtG0n5c4ougXs7ThfbPRmWMNzIhYe2oE5Y/gWrPcy9SOAFH6wBudLwUob
RsdkQxSoqIW7qS5v+5160EPNACoDB3CWyWVXIvmMd+R6rOITPi09QozHPO2VSPrBsA1WYHmoSQTX
u4ZvOmbjukebcB+jrlL8aldaZMjLVk+oBIjQU80Gzcgdg/ei5MtxS+62VcEB8xuw2k05O5og4+Jo
P/PUYWipUb+jRH+PrFrIY716q81nyils19z20KSnd4trD10r24axbPz5Xc8AD33OZfVd/qJAJJyv
9XWCp7E5lKJ8bi92CqTE4dp6LhYs8CQb4fXvBWszYZbz785XBme3BV7JbRmvbHO0syUK4zxBlVkH
CJEgqkFuI7jecL3TBNdvWXxr1s66ITdS13xSzLVdvY4HbgIC6Dc36JV98oSVcV4B2Y2iTXRocjoc
Ey51nUxMKO0Q4AS/yhZf9hjT8K7Zm9+3JaBc9SfqCtNAQ+vRz8sNBf4nfnGzFn5Gs8uuHySnlJHu
txwbIj5TWnt1d1jWMdtie29dckD7PHrXDlDU6CIbk8YVVOnww9yJhUUlpLficAfeDO3uRlUbzh0U
GlNOpddJGflUuYQ1MC8FujvX0z7s90/bikpnffW5gQPHdb8AJxnoC5raWIOXgZDXrdGn7chaiG+m
znjDDULSvnJxsFAUOlYdVETk0nwX6mn1xoEb514jqxKZjBKEHdUUMAdDn514+QVzhRdllgbu2mL0
3j+s/IBi3vA6Qo3BwWBEE2UOZQVFtxXYdUpGu9Mn8nGnlHLFVM0c9bpJ8hcCVPvhn5sspW2aHYAx
87S/62SzNNiQHCOTgsbBgN5u2y/DnsknMvPmkNdz4BkUIBelPrdqgthWsdo/x9X+JEWZNzpjIa8H
1OWc94V1syjQH78lk3uD7sLC/hMlubxBK4yhdOQoQTBzIV7Xq7rp/CuWpECIjuGT/8t5AjapyEf5
m9RMdD1agrfW0fT6hu0ZLd2U65K3ZCsWYi0d132S/Ea7C+dq9UNgjdaLoV3U7YyRCSLmixlC6fI5
SUo9DM6v1Qn2vZmSQAFmyxf1GLMOh5ZhlTQ9MbGlq7RDXy+fAissHOKelegzHN4eNMWsgDHoWUpq
K479RYmbS8zODYAeiaQ2cQ7Kk5ynb/a6B9Dn6LZUaY7qvFwqWzKZvOrCp+kK352mCuXrXjbEf7fH
uVJU/x+E3hAZKoe+SnrrQs3amSPDhkwtH+dMYa+4aoJNc8Pwe6aD3QjGtwVUUjOJ6vKziQ2CnxpO
F351jvNy+yQTqqbYLzNcNjcMjLLqjHK164wZBDF69QKvdqaevh2aF8abqlzXGCQtyeQkvAKkaOM1
6Q/6svxJEIwKAZXJ1Wd7Z1JPeNOIapJKR5Ta9QR6KdY4gEK/pzJFurtR9dmtnsp1+bjVGfDQGV+B
rTXaNk8kI69EXa46yIaaPebxjAOnNe/9tRU7O9qEGmNXvo6vBl/Xn/63868oTr3DdTtFILj0Gl+F
7GdnlxCqIdt0glXJVs7aWO4GgPSBynhI+r3M5q+YR6CIL511k8WLcAgfA51cCU38tDyFy8Mg4OVw
ivt06PZJ9a3xskt7np1pEeAnh2nR04JkRGJMqpBJOqNviEjh4IHFcLeekXYNgScmPxrZRYqL4qb5
xFumG0/Xuim1LdZHKFb10L+aD3rZbFumk9xGnLRGWzxc6k+VESWo17YCwNlRDT0O4HM01joVn1kc
Ko6iK+7I1wOKI1P6B7VuAGLfAytQhoyEpCDVDbGBZgaCnrTwnLpCvu+xf6+Q0llwE9CeQoN1sWFy
kdshOU6cludUYfc86yDUKAbnpY3F2TiH5CbhaCVc8sHtvi4OJSJTEicoi+zUNTYvQsbNLzImr6bM
MAXYQLHMfbyKbs/5LU42GsseH/jsvcN25w1ol2RCTERPP03G+XvywwOQI+VguqcSGu9yuZIpczw8
5Z6HVtBY+qiYuJkD4RZ65TWZx7ifo2Z8i28rmppF8Gkm4jNIBDhD588jMma4fizhpPYL61/+Ybsj
sd2JOr18BNmZGdKlz/Wvyv3WFfwsaHolttahKBVdcgUFGXj0s1zCfpf+1TFjYZw6D1Qq6n7PosY0
icCsKKvwcT+AmpVsFLDwreK2fHBsZixQnTTl8495Z3J7krtpnPCNDXCxjpy1XAHAoDjL6DMHlwnP
Ee02K4qewsubXiCSfyvhvOJeZuHQ+8nSNfidP0IhyeLjThiRbAT1Mo4fOeZx26gXnBK9Fk9mb4F8
NtTu33NOZt6ElnH6rcBwBDvMLsKSIzoYeI85BKh3eMNE+KXrC3QB23+mJElMTVvpeBxdXV16gg+L
V3c/L5CGUfKXr8gux8PTHE3HAlwL45PdljO6e+G5MuyRl9ZIshPTRQKXM3HH4GeoCr7aHgxNTggq
elcnQksyOlDZ95cVAvkKCV6H9vvzlL5kJiWbmha8+0ML5SAE4386fxlztkrEdm2K69+qEBwaawhe
FYyBcISmzdBFTAFl8Ci4+LiONo/Ev3/YQzI/BTyesVR1rTjiG/bLNsZM+jI2zV5z7GZ4+wRwSofR
eyJ26YMNwd0ygVNrwaeMFdUN1fQAUW9JlpdhkFEcWUgLoNdHwf4SE07TQ5TiraI1TGeYZKIIb3HN
QQSzL8kSBGI7gRrkHmyyrocA5Kw66UQPBK+yTCeTOn98WGi83y5V5XAuLdNiEw1IV+hO+KfcEpA3
zsADQRgJxqVyuBp86yy+xS18hunkt34DvQI/sTvsy8jaoA/+h5rITbvkdOKGlDszyh0eXgjd96vL
yvOxcgU9eStTN51AbV1pJrLcQKHSLIcQ2RLgef524myATTf42sL+F/I9xX7TyP5O9MgWgwcxiIuq
DbQPAIKcYYQ+hbglCITl2sMAG1LZvUf9dhmbyJTes/VhUZxS5w/gZubh2titNqrblHazAbmBRwY8
4AUOC1eVpzU2A5jC1H56Nn5FytjZqHA/Bs+16ZJsCWWJ2DKLerkTSHq1PpNH7/oqdZXDcXplFYjW
VOwS58bEEHViMsMBGLSWbrshXgYa2n+DKO9Q1LWFB6v4vzZiIkzdFqMAE797X4iBjTOPmNynOS7i
WcvXrSm7JECqUQzkXRnknzCnvcLaHJJepc0l3B2ONYv6yIJiNEtSkrGcR6bzJRy9C+5ZUzqF7ZlY
WMEL93cQ5Om3a0ijD6OhPC+KK1MMaoIh6bXcPq5XTrCFPo035l2YN7uc7AnUeuzi+GbD5tDNqKkx
QLXHSnlVe/VH1Bjup6T7n9sb/Tk8+u+cT1fbIGbS7ESaKXtLiU2EHet5giHnOz38DlX54u/eRCVi
n5g0XAnzWyLrNtj3Kc3Wdgt568uhvLKKez7nw09+fj74PRp59XTrDMtaydhu2FBKpuH5v6K8D3w0
R5k5Tm1zG//vmejoLCLjXrMV7VLoWnHR3McBm3a0PrgagbFxO6ESAEyg0CKumLvYssQFgm5NkWkM
3te3EspX2idBZm6iyex/rSKzVAqvfoSdTqBdf/kBC0aFpGcoCSai16eH5zIfLh7rgos26rbXfIT/
L0sbAyHC3mzLXxDeVDQMiqPZgir/I/wil6lYkKH5iTmq+FFvYCHAGfYTd+jkLupx3hww9nwNNHnf
6za8x/5NzjG05T1EdpL1yWuAbBirMDzAKHD85f4zMsOV7gg02IG6uVUpuHltm5EmIbeWGmL8pNge
MZGadpr1zzbPbAQAtTjVSa2jW9HCvYuqfdciRCDCYMhHCXFrzRnBdVnwZgpMboRJs5KwNh6oIWqM
3QnJm1dYc6Ok3PJE9Wr96GUB6Z8/9uH7L7CUPjzHa5B+AonXs6TCIp03nAGoFgiPFkG69wS1BD/3
LCQxDQjfv7aZ/btLUXYYWaIIWY31/od6+bqn+3LNwEJ0ki9E3eWqiyHA045UuKcrfBvoSzKryDtq
52bUGOhEXPVERL006lB23Dg/G/ArnpGfYfiWU505hlzezR9yJ0MjslMtjuRjsZaR99mqjNnJdx0r
2/7AAh5kc2XjiKMsq//X5hXgyIu9eZE0Vrmp4SIFMds6eGrUd8Ofs9kjnNQwPYaqRQcV703mCAJB
cblAkOBlIxeTEXMTQ60bT50wqdYwvbbaZNIfjFT0kgAiR7og9jjpuS0FgpN/eAEwszaQ0GzUpSgV
Bwsh/G3zWuG2vKLgTS5dwHo462h2vQK7yfc4r4uoOwZWhIqZZ9fvE9UCiDVU28Kmq6BSmY9W6ciJ
CbV0Mtu0BMuaOhOCmXkqAFP+f4+jGorwW3hapfZDYvo6samcdknlAmebaBhsXJT0vFhV8Boj+kN3
NwVjsp8/no6fd5wRQkyNJgscDEshdUrWP3u1Dy5LOfyWQYtavk2O1VVHD66YnTdWCXyMCypAfcd/
z/9yDsXvCG+FOUk20TBGUqno/0W1awWVv8WlkJXNqhkakBj0ZKh1XtSgnnXUMmXNShuk68Lq6lXT
myYXlpTRQJdr3IFgIi2vL7/RJMwTH2I8JaR4mU/PjJF0PwrZGBzuclsWF+lc/yh2lxNekt2ZlCxH
KRp40PDD4rkCIw20CJ9iQV/NX02tqteAY048u5qBpIxEUPMcs09Vfi7dHgc0jCD3PfKZos9kpPsL
YEeFElOPFi5UkzQ7SF3+5lhBTkU5E/yPEULSlAt15DAi7XvMj9LUe8QCzRNIDaW+RX8jrrscRnQW
dPisgzjfCadHsG79TMOo7tLCtZCk9V0gcOVnVWH2XnNiKBY8C3aduV7WyuUPi4IcvVaKJco2k8gg
Z7/kSvbUf0OBWL3INYG8oPeXEuimIGcuE6ywJ0Uf/BAGmrKyQevmYB3Zv9dazeLWsOBOsymJ7dZI
vdXpgr7TC2j3O7xtD87n3VjFAYZWCXSCYU3rvqcZVIXxh9WJFkSRNPuCRXZlzEMsqHqgcQQq7lV3
d7ZGXWjaeaxrMV3dKJMRROMUhJakNMbxrwWezghYNpkx+ZLCwtIdTJL/XACDWOxA7XXQRa4DjgiT
zTkQjCifAM4B3i5KahC3eu35vCYRCIwY8NCGw/pa+wXn+HnyrhMWyfEgPT2Ej2EL/WRxwLNpXIgE
VU+OZqPhrHIwlWln7BXBHvCrvbbUH44C9JB1706U2mi9w1S/ihxkHMlXSRsjU1+tRDrD9GkmY7wD
KKtcFed5U4p3lSQshSZlO5P9gkbrQb5H+qju4BiwtOj15UwNSObL9GtSoXaZ0BuK0fkliYZ0C949
uBdrZye+guMxRFT/F4TevpEsWgBsomyhnAVxAtMEHMIPG5rX5tiUlkp6QfMz/p644UDZpIxSGfAR
WzJgb1Q2xYiDLZzohai6O99HBY1dT6J4MGKaDBWVAgc01IkGCpwWMSJfziOb6SBYj1NySkJHZ9dj
SkWocWVo6+26SZdqIusFKz1xr2h37xL/4/CgrITgpTfatasac6IO1/qep6sbWf/i9kFQ+TZT/aNe
TzkcqOFXor78HYqUDezTJrdZi0O8736+lOOExllCbmeMdGOZhxLh8aZJ03rdSafFi6ZG1jITlgw8
53hU80W3T+FE0TqZu0f1UGbr8S6FkHJFGbIWq/XJp6F5rcNk4UmTUcMqPcKpsXUBR6OA2fiXA2TL
1TJG/elOrCQlqj4D6sWAsf40OMZs7YWG/9qltRq7ZTmRim4FinnQ2SLfu6ahd6/vzYA6V9550R1B
2QtOKimn5RIC9a51yCVzZxDBhrT6dUTRnnQgy5GZjEg6WijzP6csVsQ5+uYvXZv3wvq+6GoB9dQZ
nvaROYySKSsCMxgt/C/QUK4nGRJlb84MmKUtmixOqd6jbkWOgII7PEa45p37pTV3oFCpiuoF8nne
AQxNRl+q43aH5ftyUDFhZYs0XsR4RzJjv0EpA/hrz8D2Imlmhac5WLr1Z3NmwvE5d9Jgq+Jk4Gcm
qFP5Txv8wkdJYRNR4OzMeMsroACmVyqAn9k5LvJCIe0M1Tvbl40azMydmCCVbqJ7zSrVu8EtpaeL
WVNjaTqmmkwHfhocQiz03dFxx15xM+dGFlvcqHo9bTS2KmPP84+AVtknA8LQ1vaxoz2/ZRAPFDex
WHjOi7YUeA0s10MVoAHZsjowOlX0h8fnMn8WcwpSkQ/d5HSI+HZT54PEFyZhMHRy/r25xrdq2dPX
zjZk2a9LSiZH8IS8q/xxVqc0jSkCPZaJT4v2QLu0MqGWAhts9UkX3sL7qRpI0MPoB+kxGIBNoSRt
qObq1M4xbaIYO/ObS2hqYipo0O06mzNpuRvNHqc8ML9P7ETSv24gdrWTMljeeTcQHSgCH17CTMy0
aWrYIb9xM36JWdHYFhAGcfUOGzkKzCd3elzmw+6oDIxvKp4iev+IHSbcNH1yKQAGe1FL03wFDztn
ttYiCuPBOS14fMoeuEu3H3hZo163zjEMSbKKXd6qdWhuOBsR8n/VzY1pCLIroeuYAO3o3Bu0xFkN
WCxV0EJmCZSV98gb/DkY/yYbj/BdyB3vfVbmU5NmHGrtoV7dz+DPUfnfDMWVSJ9kDRNNLW4Lhikr
aRx+WXwbcfcqEk8CKE/pMfUo1SQnbyYlPhzyroxbm04Ts2BHUnzRYDJm7O8mO+W81lm/BbA6SYnN
wMxM/ACyGvs5pTgL6jj7drqBllbpUWOyfuYR2Agweeyxk/wGd2um5VzKF0uLruv1nmOgJInt2I0W
N9HmkuhJuLE7cmbV6G6umt0bWbMcpQz669de8ADh9cgJJ0V88BOIeGqFSQXzcUWnLCTbhs7zS8ZL
e+1CcJjG8n/6PY4Reg/OMN3wKmasnk/d+Svg0Ln8BNypIK0EFXk4ekIpyOp0RGhs9XwDUoP5foUj
DzO1LTsIdEPWd6QjpvbW5XP3Qogm1jrcZymacGYhgg7Lr2EW3+G1RWtSGFUQ9owvFjCmtGBuwNpD
3ADmcgUC5cxLAP+0BWhFXtHa1i2M44tiy/GQZOCODem1zPmG/GO5vDnqxoxT80xJukxSC0ZuvPfa
yoI4KdxeGUnH3qi4NQ8iouv9OkVmVgh/4x6VwZpkQtM4R4n6wVnKellpTXNP2b8rtvex50yvpgDw
ifj4d+tuAEGqBfPe7Nf6/cGs5Kkn629KcD1iRMdnpfnBEJLWk2Uo1MWbF6aht5vGI31yl8IyX71K
WvfbGWguvIO+63biYaQQxOHDWu/IT1YprcFNbI52VHYyQImzS1S4AHOo0oCuTpA/+zDmne8v67dH
+kN5DOryVgUaX2yQlwFikRsSI7pOrB/tptUwUMTbt6e7gOQ6fxHYcKG0bxbK3Ui9NhLUwPyc9c4c
hWC4TyZHt9k0Wnx2Yqj0YH9FT4AlnDOdNq1/dOSd1I1LtdEtY+muykO+LTagPWZJiVD7rVFb/iJE
+x7OM+dB1GlO5WlYg6uqWtrwgRtyK3DIXzrntCHDvUopCxrd9SivvwJ+4r03amoauvK2ml3xYrch
/Gdg1yXhhvroaXMYdH7LR2rGwPkG7wfjmDB3jtUYTtk/db8+w1oC3UsxiFtJsHTXj/vQ+8RZyJWU
WEs5uWFCU0w1mvHDgdgfPNlfPfzfpdXkqLRxOvxjtUxFEeAd7qcfPHPUwItdClKLzgYU/my4DTK2
OhlqkeRcDeXd+GmTc9TiQnhdBFYPXjyZgGuAHiaEm+Dui7l3LC9CgUfDnwy/rJPkLvb2yn9CRKfB
U1fzhJGgQQU+Qggm4/VYMMJf2dtCrAjhiRgG7y2xya5iwBaM0NZ0VKxUeEovJS7kjOaGIj99BlHP
VJHlpaCUDqFtGWSluQbdJ4dkGCX6Z7Bwspx1LpmYoGQZgz4B2JAUKucX8IgXM6riVsqb4VFvwy7Z
VkgfOQdmmG585yJ5k4210RDbn1C+mc+cpVPaoF2hiZ7Xdpum/CwlUpXOZyJXQ2eMgV3bOMsj622k
cC/sEcrznW5io64JGt/sRbNpCbx2nERVFm8kOW89QYMF5SqJQNmC5ZFYxu3brfiUfOZ6ZQYNRynC
E+G6PYiMFwBMiB+2+yKv6L99Uoi04GHchQHE0NFlQ1K8491skBvh2RMWm4oMThsJNrMmBv+ZDCnS
hEYnELlGvFfUT21efZcXiTob0N3rwsK9VXk+IdmyDV0538NLpdWYntf84nuc7qgiHch1GrhEXYwr
Q6acu5tJft+h4mruvF+Vw7avBGodbfbDbzjEKfv8gXTy3rYO64rBMl3cIK6JUCBbLGaAw2eouSU8
Ux4L/R8B0S4OwhN9bU6YlSEMiuFQ2YUswSgVBzNal6TwX0rSQWVteca+HQQTBtWlsTLjgN/lUQjj
ISgAu+wCLvZLI+ZwRcoUGCS/gLY3ZBVIUlmeUEP7qEV/UTS/aIrxTrUv6xf4j9E7w1Af+jYQmrPZ
dZRt2sIYutE2WpTvPj2g6ROODbVOFzmL4q6qzXtQBnXBU+JG8ElQWpJcGsDZ6bV9GGDMX/NmJtbG
iyYtIpL2BvxhyURlyykfXAKNhwCLSMz/Iyo6qLh6cHJuXIedshWYaDKJzV4jdRwqXwZzrguG1ZUU
8f15RF1nN/ebYfjajknyv08yzpqqDpdc12z8xL/Go9kniBZWMdjXVr0Rps+LpdFmXBYH283K1kuU
Iw6SPo2CwWKFHExZ8NffvrS0B2s0En1gIJ8bius6dxSHmO7GLe8hZya5CR5lP1WAnXqBbnRLQXP5
M8pDtBXfnjn2SQ1XtckQeamRUlEdq6kF0uqCXN3iLxrrXTsJw/IuYhfqAK0M/wJuG2nMSvb+YCSh
beeyvf1aZN4QCYAWITfC10snI4cJIR79gEw+u0rnZBbpnAH6/SjzI+T9m3YNfgM74/lev2y5sXAF
GOOGZhhbaqLoeDGCYwYqqR6rliu7S0E5v4rOv44jsJrOcfONyZ0nhiGwZfjuogHOLm2RCFbZfTgu
ef3+oznagaLH3IH+2TT/beXaCV51CgQawfE64vbcieC0VS8fNuMes4brLwuISBLgVkKhhz8hSN+K
wieHQDO1OP0pZxhVgkB+iZTj2Bj9rBxK8wFLF3vmiDxQq1aeNzPEb5sqFbt9R9w4KZU47DZ7tvgw
nTVgwSP9I6fGGbCyyk3lvzDDJYqOhb7bGGgySYaqKKbhuoQSWxF/53RhlvmBfteCSlc+MHsXhsg+
p5b5dAu+SQLkjbbt6Zk7n0+NayYe2NW4awORr+Xrx74O5vV0ciyZvzqGgN7TGy+ZvZIySFEk09bc
W7Ol4/laWOpGy5aqD5hd/kh+AN+NMBMRxifKizMLifn6seJnVXXFI47wUYlmVku5TpDNjeUQQXDR
kwPviCGR9UfnaRiz8tj3/u5wWySzNB6jrfgDvcSB+fQZIVUArPsAHZ+YsULbTw65HpXHxvWQ+Hx1
djOmeNzpo53mH6FSY18cibzqeMa7Mg1fXsKw5GnPJX58+NuI+NKy5cQ6FNa5rtkCmeG80ufoQmVG
+n03gv+8FRlO3dhblZdG8NrRfGAwVc2SSe/TbznLRzkZPIZBWSIUglZ68II0jR6M4Kg317RstM7U
oPXe7kAatPQXY69S3fUgmt/WLPU5kIsD6X/WhapMBcMUP5vijQtQMy3kPOmI42RSb7HcS3JOfOEV
vGHzcDoFJoQsi96eYLU2lsz7o5B4GPSD04+7DuYi0qzxE2y7+29Le66jXx6w+kRDWIJe8cYADlR8
COh4BppJBvuopMfZtjcB4afCTpEKv+ZGGP5lEDh0xFkTlvZyGN9n1AVFWF59gbj6F7kRQnnL1gPi
EucfwslBHT+QIc9J2hhffok9B4zxsxUPZLqJRttLgfzhYly3bltwI+jopqPnilcjC7vze+Zx5wZh
Txt0A1bsss2OA20GdpRnQoqiobng83CEaMMVPHKD8cFY5kCKlEZOm6HQifXZY4VTQaAAz+gsfH35
zBTNLzuqVYbYO9PBJvwl2DIizgMlN1+0LK3TdPEEMujZ0FXzGluOf3POyTfXwAw9dxkSCsOArupL
0zK3UtpUM0X+oxCleuUbowMVoWsTE3u1ajfj+NpXR9oWRIAS8j2+jEV4607oXdLtLLItk9Gmrau3
Fbv2TKO2hQPFUnSJwPuRBaCTylLGxMu0r92fYzp61s8BNofg1AVz3O+im3UurNFFfjI1/tY0xbgT
I8qVB04xvkkMqBKT6XgaC0snZOAXtx517wK5grxytsfaTMEgSghbbzI6f0qqcW0o6CMHJPokb/qb
IzaDqT67lg62kxW9llLDyYyXJJ0V7Cyl0HmKZYKTsfRhse8HeyVBbGl7yXZ/wdi6r/sKUmhfv5I4
DSQCZF5ikW6WuJMSe0Vw7/MQFvq7dT/aEGaQZe+w0U0S3YIet+YU0WMGzuAPC2xk8UD695vM/YvF
to2WtJMK/MrQNDOmt+58JfArrqbXGv1Y51wrZ+DXEPL8Xmjtox0OcEb8zieZRh4vKMdf16nQFmgD
ncUSMtGL75G2Xs0v78y2tD+rK+Iki/df7LG+N7EcDU0GqcX8jABO6/SWNESw/cvoTdC147l+6cpk
3kVjZQWmzN1ti46pT+B1aRVjuLtCcPfOgRiFl29fvIcrQLxTfTBxcXsRMT7sBg0iK0WqZWYd4j5K
hjB/La1n1G1CMKavyH1Kkkp58d84IbABSnEvEYQHQVj2/fX2V2kBougI+1yaPFK/vOGlDfxdKkdT
4NYgcPEdY4e3KNaf0zImwzCZWKuLroIdkyZZOrpQKJkz0niFAv/qBC4G9+XkpY02P3aAFLJZO0ZP
nZcRHuA8xoLwV3ZbKPmWDEq/HiiWcLlwMnCTnNWBK6WSiy1lv1jnkZMg+xXmM8EM3nFGYN7UD22Y
rPcfvUhX9XY5GwyYu/LDVdBS2Agk7ILisZNr0vtM2TREpZTjA1ajG1Iq2Xmud19QmDxZuUH/zyTE
nHdQ3yXHLHHcVjL1wROTU/h0iQ5SRipyQfJFnhIN77clZDIV/3AXCcsyEzAr+Q6VSwQEGZLpvRxF
Sm5U6AusOtBcsv7UVR6U1cyym0AHZQz4CzhICrguEomw+xG/yL8YK9aDv0nLBuO/K76HZVlikcmE
PRtzS46rEFD4sO/raiX3TRshl0qoVV5LJieGizqb2Zt7K5YUqNNfbTXCLJcgR+2e4Q1bvvKgf8w9
okaR/bumggrX7LaztwfkF9VPCuPp13mZVlB7hXJ3eBj0Vte4CR2NOdEGDFAIupn31Gf2rsoV4AFl
eDG+Jnw/Qir+f69lGpaL0LKYLLHU9xyHNMpde0tm1pnFEv7n+Be4K447/oDOIYNs/p7OsFHTvt7P
FYTtM9XTQNHZAm0HFhq9mdCYbGIp01t7Yhs1pgZXwtHPdBbBoWHrSAKr/cBZqLg7we5mP3tMZcMu
7k10tEJ+/L8J3yGdAONSPx9DimViK9a2iKTUzmnIh32OfOMpsZJZbmREdXZ96c7PB5nwykjx2EDG
CEKx2+rKRP8pcNnmDdA3AwOQSvV+KdaMEL1sCbsT77UYwZDeIIhR5Lo/EljbtkbH4iQOWW/bWvY/
cCay925VfNO5sC64A49mK22on8XBvd/+3YFlUwm8qZI6JXErrk+TJvHNejH5dxGAyHyNtd9DQIbk
AWOPfZVgdR/Ju8C8eOtTaUfoUN4Ol14bOH1tywXOqK1FQIOoO2xqgtm4m3oWpUa9MkCOfYe+RsqK
je1h/j36mS0yna60Vmfr6d5kdbi59B6cNITbgiifvLHjgq/b9uMLkjMQAM2mBmZHrK3Jua1agft7
YCmkI85ArYsY3PpQbEQIOBzJ3aj216dN0mHBssV2RP/ydaOgMFW/Jtxkvx5xxqwnu4E5OPFfLAqr
Z2Npr4pA/yj9RQV1SfDhPqRrSz8nXN4/Z1otrQGqz0HAb9WvEgTYIZbMl/DB/HGdbKYmMrnCMZIi
83hKRgqCl/dCG2/22nTQjIlftwmXvdhdYG9y951fC2hcpWo8hoeRnoqGqzcIqrqHoPmbMh8Fl6dN
NwbcHQcxr1rMBrIiHAISy5rPc81qYFLZsz25Q70bUyg7Tkz/LGaG/QyjD3o3ujo0gXkBVSkMDF/x
1GiqgR6eQzqkdVBy/wLiXETfObTIJlZ7eRZxJP0ZQv72hOTPSBLKOCRLcZANIi9kNBcsncp9elc6
pP2bf96NMFULTjvAHzARE54yI3f0PZYNq9hmfOO7lx1TdlRbLxUqegs4MeHQpvjjDdZPcK04Gjw6
p5e0SUWfFpGxYWMeVg1Oaq5+D/t9FnsIlKNbT66IEQYfd8W2fCXxM7ZuJD96xUsy9Oc9EBcGxDXr
dE5fCHigEcS9oX3Jx7WFDtYkuGOeon58q7FDuLmdBjLXvPeaGgtXSXT4k4len7Kg0YeNKnYo0XYC
3RzlNBHAEZw0xqiERdK+jXQ1nv9BzzHzd4tRL90SLBpCqUIuUclZq7dZH6iAb16XLiTUASxMbe46
WWPaI0lnL1WRXSmxRXFWmtQPGvBlIuXbMi/LsFysWdIKBXX+ZzjSbRKYIK/SmRIuaKB1tQA46yju
S0Tb2yndPzK6cUtpjrha+nv1NsW+ogb3Sy0vpIdmTK5naIACL4hcs3+hQuy9gkQjLHVfdHDKs+1Q
+P0ZoaHZiL+eVL96iRzO3ltxQde2YOEJd1zUPpvfBGZ1JRsLYYiJXLbJZsh7bvFgbazvS+l9R0BF
mY32VDiv9JqEV9HjNZbpPtnHfbt8RC6ms9uulPFBwCIDx1nvYgGFie35GnTlmXwKfxlebIDwNcjw
mHdDX99x6Zq9SCS9TjKUgRtkLIEBy2IloCtkcMl9WsMyDohN64TdAD6J2Q43IJi2ysLktPiMqaJv
4e6NW8SEIur4WnFS4kc9wuxEbQVYZWgAw9srOt2hVUEPzkdiM/3Gy7RhkaVP8XNy0zJTDiSpBM65
or2yVEQRCDKR7a/YyAqby7exd0Snt2K9S7+LNJ6izqG8qQ3f10oRiJSWktHzyK2vnfK2dVcvYvSD
c0tcFc4Pmwts82mG9POsb+OrbLUQyC2H27dguYKU1DT5gg7joinF4ypJhC65ABSX925YkvicKl81
1cqDWIHGNfLUHyFzfkSj10mUoeUItGC8XkJ1ShHqSuRYYv6cOIYcL+pJ+KdtUzdV5WI7GgDTPtr+
2ThyL3qiRek+IV3Cdk4pCVnveNI2BhRkrBxSTlgGcn/2bhb5Y3l8JNsQqizeCXaGsIQYy56rRi4f
XVyXO2oPLfiiqIEkzTuCj35vV/hB37MAEVK1j9pU3ZQfhtGsT/uvLdFI5qpdM9OPEaYvQBLds8bm
//wApXXiMVMVmvUA/qiPB0/kC/s3AKDvM2nbDHTbMD4Bisbh4A4/3qwjvGDa/laO2S32HkbgzFY7
hJuNrcuczwz26JJWa9iefa90FyjmMQbmhKKe7gIJ3hab8tmrQIXDMeEYkDAJwfCfA3H0vJ3ePwus
Yjwwnt+fkmHgvIW70kzWA/feRqQi8BO4TOljeS1KuwHlGa51/gNJf+Ii3jh6VlDLQRFf7VGg6X+0
6nEqNdrzIxDlsMB8cASjL/y98l51eEl3zjtpLaUswxDaCQu7OHEGsB228TFH3tj4dSmO4yDUH+QL
CUhDqJT6CWKWjQcRs5RDnhhWX8Jgto/lfhtwIDzOI+3tX+KaC4hVWfKfUoRvbCaSeBP9Qqtif/Yq
Q0ulAAMSOUkr63500N7zkuGnwrTVY9GxC7zOdvPEn9du5uMqKfS2eg2gH7BHvarS9YjNN3yWsdAr
Ho/tx3icabG8N/8QstpeUEO1UciD1/B529cMhDcYaHefwqCRK1WkmogbDF5En05p5hxE2PH4oaXo
xzqrxiRiZDo0VEEnk9hyuiRyZA0WB30kiBCrYeU0gS+mxTULMtbk47i/r6TKgRELd7jNe2kGK968
R7D9tsfZOzgUol4X6Uo9DYQNsOm5hb8E1youNIy/jkYpMUQEkEQWz/y6G34dkgOY2VnbZGGpHHB5
xigN3MkZ/jHmptPCGCIbNZXCS6VKR5fVf4r7zKiJKR9x3cbpjf39K0cAwD4ihjvdvFftm9DdZ75N
8z5l+CklukpsrNyJ9w6sBkAtq8+XjUZIZcl/A53zY9H9MP7JomPgQ4MVVMpGfJFqTmcGg51Fl4S2
mzB8GLG6Jdqvx7RkKlV2UsQGOKs4wEsZ94gu/GrnGwduOmdUUTL2/5m7c6PJGpuPxQxg94BLXPIn
iGDREaCIlEuOiKfSfycPCol3CYUCTURCTjUYkIPdLJEnX8pqP2pzMDZQF7qDEKaEkwxvCTLpuYT1
+K41MMK1zCfkSsLH9amd7iYMBG7JZX7wUX0ePb4AJJ5RTMmtoaXWOSc0+UvggNj/OrtCTqpoHP5m
oPBsYFuDAfa6acS3HRaQ3+E+HNSSCg6+p4YGvsk5Cy40QPz+ybqYuHDj83o95Z3fEJ4aukpUIh8z
vUiyRpCKMnxUHqwX7rAF4VwAv2Eo2Xif7tYtTK4F3ezZ2hiPHeWTkTNbDO2Vo2haWE+XdDqX5zBO
7BNNNNNCQntedDhm57pPHfc67Vh4ELHQvm5GXOF08xtpjvF+Tfz6825nA7HJxrBjK3e3tforX8T2
fTJLxmjpM2IgT8uCnD5FZHzQk03h/i6rkBCMFT8Q736JaflwmPKZQrM3PvaYSlzrzJVjBzJhpQGD
v5Krqp0A9qzuzohBmPY/oB9ALzESuRAYsn67oU6pW1c9L2sjj8gmC5jmBYayTtnDmeROAN6P6vD8
AapcN82BkqFHIBNsc9v7xodsN1aINqbY/GT5esnU7y55c2WDSH0yVsAF3N4VFDdDIS0M71Obbota
/+UMVqnejw9esXOceDhfL43LfDr3fZvaMtEFj4FMOy4+rpPlLuWqIV44vkkz5LXE/k2MQZMI6wDr
fvm+tBOJaj1kzvpUqoj1eSGpCvnof6Jbrw1J9Lcd2gkmYOHO8wMOb/b3qwe+Tl9yxREB/95It/7E
vuRIQCurLUEbfSK6Nr/Kxv4fsdDnIs7E+v3O2VChbNeSY6cd8cceaLTLkxEn3YDFasBy4OVrnYF+
ykWYbvyC8iz3axUGSq4aGrFSMZ8l5bY0mFqO2ntRV64WQg7JbiJIy+v5TyY7VO3ycj6dHng20WyO
FTJcxZis9nB4IlfUTv7BJMe8SrGHfPvsYTAdrIj/69oUxfFHnolX/0OEATE5c32n5LGnJGNfgIi3
y0rujqrvXx72wYYdDYcFSY+7qm1ELSxm+TqyHMXOLILU06Lz3Jn0p0lVZfdVAa2xrklwQU4ZUs0A
X0SH0tbwlPKQR173FVcEd0dh2EwotZ/JuqZ8YsPmNHa6Dkk/rPhR5E/m1CqX+WJGF4ph74AvBLoc
43I9OsohXp6A4tzSuJoTZyBNg+rBnvyMl0DEjjeTUIHPdGVC5i4kfWQOfjO8eUDUiX1hv+8AAXbt
nTgB2DBl86HmH1HnyVy/pZXA41/kIkHPol2MQ9hz12J4GqBIHB4XQ+pCEYn8qUWsJPHXkmHxEihY
IkT/X4GQzTEVWQoYDlm4cqz62CT98Upc9uLjE/B4VRdPlSKAoMDhJZBCsJ1YoeUPZr1FOGnPXv94
IScskaGpef9b6meTLYiUOJK6l0jgsOR1+d7JonJJoti0JZct0YkkKI7TowjoAFLctgmYrhXJk5vE
NGbGP+jzV/sPlQNqjnHDwek0jF2aGDvjwLshKmMNT6x0xxirepkYR6w3wLccdyL43S1EMxMQOyWm
gtFucxL5SCDOBsR0xQqQ4b376qTQQT1ltFfzsyNSNcI/QOykCTURNl2/8DKpS/wFFeNwe2B7/NS3
0wvYGGmODdsuU/d0Po0ZPC9ky8F5A8p8VMJ0fZ/Q3ZvwsxX0sJ4JJEfJ3Gl+CSSkjblMJJpXs3p5
jArZfHFEeKmNES8YPRosLMAVAtN0sw5vn4Dhe1Gu9DICRjT8qmiKvSYfT4G9OVFARqIKpRI8tnNf
vRCiNUO/zn/Wy+TPsGSW/HbobKG1cfecqFf/qDvIP7q3YgavX6pbBdNE5bsopxbJu/4tS4cCMa4o
w4ScAWT7I0zz7ADhVKmnkoyfgOg5Vx1e7B008vOhyrez9HV0+o+Qat2xtTOKXLE3dsgt4cFuFqlE
S39yAUtk87FME3ZHFIdsmgEFNQeZQjh2JlQJSvGd2s7YoVAQaP7n1KkT6ujPh78Vpok9iCfCZU6B
Ajh3ibp9mTOiAWo998tEVt8Tk1y0W+PXzckvpSR3nImL3udMGQKD6kUmto9M6O3sjD0EfFtP7Aq8
JMvrTQVEabZ2VWLIgefZUSzQ6xASszW7iJzv8WWyYq46tXwL19IAQiZ40hM12eDD/yPR3+rhUFp5
0Np46K8swYSvGCEA1ybE5mxHRNKMb/ySyk9RpLyI7vwanm8b+eOXJ+VIS9Sh0WKlJFlmrL0G50or
0t7Vfe8Jx5RsV42qm0Fpfp6ooTQlx/x+udCbIqLuKNOwIvynGTEyxzktcAGQ0PTDYsOkWoRELZk2
GxGgV/ys/f83EUFC6BiVIee9eQOLGVG8Ws68HshxP7bnOhUt0MQPjxCw/jBFrqCa6T1ZLEUDmB2j
2q8ESOitqtzoe8qrBzELF4DnNUyHKVLhSKrFc4Lm4JHNXxnJdd5RP6PfioW1+gqkhqGHr9cmhYU0
mfNDLUFn3lwaseczyQhYbdv91QSxLVCeFC+X/yFA89npKy3gj9c/oGKiATB9pHIYNPmZpCmBSHdV
567t3tjfJ9WmD+c2OTwg3pkeQJmfZ0e9J/veyTSJKA7d75/GTeD2aVFimHBJUSV7FtCUD2tfTRmS
LCUSt/wjZsYTQu7l7KcWQFD92OpjvLucMOnSE6eSRqzqb+5SSkutwIPVT0YT+nYTreF/OZ88wHfw
PFa3CTZ4z/6IOWlKYa3n2vWL4IWqY2/nBcKNOfgTxzSLUTj2OwTCzqkmlkieOWsl+JWf9gYpoSjx
29Ei2kmCcOkhQJSL3hgJQRCLYAZPbw/6hiY3GFJFCmVl+CczakrMgEGLElH0LCHmI/Aul9GOPN9/
I5BMj5CqIJnr62KHFA0ZePg8lNo8o3EIm7YrFJhFLZneyYncbsziUcA8H3d54S30nYCWLQdZ1soH
YW4HRgYvaDzwnhwVVZNY1GHMv9ZMXGzM3spym8P+69nKdBcpD/+nknF14N45js7n2jX7v85dWAJ4
d258/Q9g+RrejGDOCmAEQhAL/bRABx4Wpe8Asm96kip8/8vZAyGSNxpeSMCPo0Yg/Nc17F2QJMUE
krjFNie6Hl5CZMjV99vvcdWyZAWD7Y8JOob97ntzbUCzDeFG9Y6vuXnem3Ou7Tm8qvWB/brV/Q7K
sUSdmtsO8EdUvo6PuWC5WyWrLkDuVjZioF65RwipxkjAxNOuNqSdPwa2qxw9H+m8Gkp1P779l3B2
8odCSF2rgIVohyA9rNAY27SF+6SPUVw2l2sdh70cxxfN+xmA/fA5eefReEW9CsJyIIa2Jn6JEb6w
DmKIpfJKWhg68cq0xMg2fUDdPhHtZwZxA91IH9TqCfP8uQsid+/dHIb0c09uWggiGlNAV/mSc45d
wBnJoRyMwRzhzeuBGVyTswxJwpOEonImlxTI/8SJeV7wwP4MFTMQ+cIHZ/mSShizOBOPJUQjIM0i
mlGZGudwfxUrzOHQ1pdNRqh+THVH6kSSd9s/ynrNosK9wWTqWXXoh4AB3d9CrlVm8dCmG7K6ZuxS
4/qoy5W24zU+TJuF9HU4h14AYd6wTPIuujYjdVrROyHEhcFx/5UhqW5b0GgUkVvJSbxvdVcUR3x3
uYtgeTJAm8cA0tn4E3XqIL2kPWbJS0+gXE2EwcePy7IqtOSmDO3unoW9mM6MVx6vRVgOgSvw9znm
ZKXBuE5VnlgYEjfdNYDQ1YV+zJMg/QEzAfsUL+I+dFbVCSNnI/92Lep0GLsBMnt/As13Z6gYPBRj
hTjMgICXJUMhfLJDiMg1ytSY4dSJ0ffjyQ85aEv7lQ6vIgYLOENVeyoxhm6FUbOQG0am+vZsPMk1
W6DL8mTJ73pJnZq8742Sxa3iQ3SENxzH+Edg4Pbg1vEs+PrU8xbcgXYNZIFXQoOwOtkGCgmQa5ml
RMrdx8euZCEO1OmAixLYJnmu1fO8n2lqBnqUJn0OXxIsrr1GG/8iFDBxDanABsEMHXO02nMbfRAu
29EzgmNmFngzCWvP+Qz2SvHLn05TGDOo5QpnAaCVkaY9iVWv6ia/bApWceggz3Ti8I7bCZE9O6j/
x9/EoapZPdLSq2GKZGf56MYN0NBNV9PHbg1gAExqdI72i5YYJyanGQ9Psul/F1NolyfhB2V8AII1
sIqGQIczr6PydCVuO8ku1yYVDesMqnk4K1oMqipqCR8avn7xi4z6I9+IpQNlvmZqv6X/DQHa/kTc
g6/G6MtY4oNZjN1OQ1vtXmiJpIdbvpawMOFinmyxpR0MaNTSMifkg4Vh/aHPZops5IDimeMMudPv
RiDJ/4wbFE4L0fAt+vG2H0jYBeRIt8rR03Zggw9m6RbeLGRJa2m7kd3erUfsiu8JN6bLMYaVmCXS
cUcgm+ONaSCi7OBj1RXBSjHBpWCAPw6cQqMd/yGu+dTbGQvJ4zz9AYooR4Wwok3Z26yaxwi/T0EY
YwX4niRFxpFrAYfR/kTItW8Sny+GgIwlXHXDGxyXlz6kb+Gr/X04IAHEYQXFMHBBWPcu5bRWVvmX
deLeRMthzs5/A1yeYAr2Ct4rliljUxVWGOMZUM+iA6Ai+7GdS5Uc4aPZD2tvGkX5wf0qmPNFkTHt
M/u02aiAimujHViw0OKuBLvbfWnz7mL4atKC0Th1kHXf0buOArS1Buk50XmwtmgMjzVJm8Ko0BpR
b/qBhmdgVarmDlzYtXFWwpBVq37LbxYIr1PL4F9gYOg9rFUUANBGrxE/Qs33q12T4SsJhlDY6ZwV
EdkF2A0A1qIdoVj+BUMM3keagJYJ7rqd/I/GqP1daWvMMVRJ/+fGkjALKVYja0esXVrHK6Uq7EnU
vq45XTVTTbo7C7pmzYXiOBOFG2dqJDnZLOqp566TtJqi4ZHKz2sWDDfcWX/wFz+Uq23dLO3T3URH
ERP+d5tsHe8aVabq3ZLm66ysR33l7lyX2saqXf+njcgo7uX0or3ud+Fk+4+FoeJF7R6RJ2AyAI3q
A1YUZNsGA2CGO/rgZoefcN7VuwiQqoOfcoh1mbSqQt7agIp1B5aQeD8m+SqD7nNthuWsdXvVUhf7
Vn9U30IkXt9Mvu2NlOo9/CNznHnruzXNvaebZzKIoKIo/qD1k1h3KUhbB9Wvvl53jq/iSTrk5/Vb
zhupx6yvV7grigKGXqPS6IQ93OoMlKZVboFMr2G6Mtniua2vQftdeVLtBeBfvy8QN4+IlkV1lWwF
2tvw75DBnEa3zixaudQY9GZSLLDoLv4HAzlUFLSqo19w2vHjyfx2OAM9xk3YywBG32Bp+CzoXc8E
61HkmxEH7GjFbrsLya/Xki5ARmJH+r7kAseCq4P9CKgJ3uo0q8fDuDGoQrX9fZssOmZZeGmTbNEQ
WWN7nN9wZAn2g1LjQUTn37BO9q2lMJ1G1CF7wNW/yGsxgzP69gh0CEM75T61LRxazDX5OM2FFY0U
t+0n/ppid2Y5uHoHz93WsNJaXoDbfqged/Ua6+xEKwlf0VqEAlNKysdoITmIIAmTfWaZ6Ob+15Z5
SWlBv0LsmvxLVO139vMEnMqdmE3/gbDyrq/QeI8vdY3mb2rmK0JJQ23komvgNKN1c85B9hiBCrCV
KpMlj9zym+vkBjVi//vsI4BX6mi6S2Ycvlmx/xJW/CVFL3tl33qVzFxnb2pG+/LWsM1ZOzwMVzE4
ChuDnosJB3Gg0eU1jVRtnTy8MdjHvXybFK26EsTYoOUkurG6JPIxU8NNVkzs58jxfJ5CnjSzgTTh
gWAqknGipG8Or6ohw8Em63ZHnVrN1Zjmcjx+gpPrTWmhPyY1i032jce/tkA0+BIAP1JZyK0Y/dCt
GA01LImyzy/vdh4yh8a09wEpcvdB41Bas8bQUhyJwvmmjJTMs0LuDeMDOqCfcTe/wnkLP90DI1nO
tepOYfxRWpZMXlHQruW3JtIqwt5tb7mKM3/hylI66uyEtz9Gj06GQ4I9605MEUPEmRGaKMuhsKn4
cPrl+h4N0LwNiGRNq4SKoZ3JLcKglEvAFaAcNMa/N0X0d2WnV6xC6tRTlw2g1x/uA2Q7N8o7Y+O7
/lYkdliuuN11LaWQmKd+BEqAsbJjz8CyNX2pWba60XhNwut8H92+/VJ1ODpgcfhyi4xs7KuhRVHF
cnAaSdCJZgkRVESAHLGrRKDLaAz18tWYZFCRAXSOqvV+vQeOZu5bu/jCn7QwK7Il+vN/iLmAbrGx
YhZTZB3eAcgtjsvWwc7h4gV/vQB7jakV+GO2XDN+G6OEQWZX9VRPYE2SboMojHfdxYVaelNeOsZX
0QcugjsF4w3u4AZOVSSIQkRyWzeiRXnJ/PHkkAL3QHcj+YXG4do3WxPxBGaKW5rajK5gbHv1spON
3uOZj5/xUj65VX5xDJ8V3/A1GHCAI7a83HxHszvgyr7kQ3Vu78q9ouF8nM0+O2myIBkbxftlA04T
6KDkizAeDRjiIqPgjo4lAZKhYux5hk5cwwkc0hD9yxNJcrEMcwfBWb4rQA9S8M2zDebYdJEJAfkB
rGHXlOqQRvMclU2VLyTcki53tjEG1D9KXXIX9YXRK/KMm9li3LeY2AIiKR9evM8w1tJLi9PEZH1d
FADYokaPOdfcLOurEXvgk7izJnacYkVgaWvDshjgeTi8bz6OMT1lzp8gwBRASOLX8RhZUtGWWLht
4CRqTCC+ByCKHinZ27Wmy88o2/wIElc9IuEYDxQa1KDEVSSVw9zBW/u5pXG+1XYZd6aTS6CUdWOG
Woty79DMLFUeI7WlDQs8ZU5usby7T3qVx9/SmGVj2a1HAbwdGDuRhYqJ4QQYBK6CD89dRtKf2TBm
S788m0aazg+scYGnfQDOL6SmaFqIZUlfIPFtKvEk9geB89mvS/YCypu03alD5aouB3J0Joy27yC6
xnxXBzG28z3iwG/wti9XzOWL7G+/PU+uA1vD3JOKuS0VSrjgzMDF6094xvVKsYix8GPHuhCA0Re4
lWd0HtHfwuyHnz1/CuU7pdehhAAOVoGqnsFCbyFVNpS/E/mXQzUNVEQNGqyxVYGv5wTmyAYkXFNy
1fPzP6t93FQ10csJzT+wYZblCt/iJUnOpLfr8qzsdMWxXYq2i5Eox4oepjzpL1kQmvuPhFOawyL5
SbvCFMbJ8pZ1+4Wpwie3emf+9Qz+4jZ5evDaOReoD1O8E4Bl1CsTD5bTOllJ/8v+KRHzNg1pA0NL
wqjDQEs8cvbbIAr/z6PXTpMDyNgpI65v9/MuTy3r2SEf56WqaUlfHtqUFKSQHrn1EjCBtVAoHMbG
gsxWKheaYK0O6P3cCrjEYQTxHIuIDbPC6uRydLWY6m6saV7C5KWAuR2shF0sFXCkRX1+ZT6trYnF
ABNhRGMTSwzB9yAwtEOSVfkyT3Y12AwKMI5Qv6v9SukbpE4KOuh0c3omb91daLpXVsrTh9z5lUMT
OXzp10zkTF9y/H6yNkh8Rt4QkzFSyPdpBqcwtaHddWC3Qc1flbi4L70TjpU4Kk+qXfUXbTsztbqJ
g2AHTtgTIJGiRfzqevSlZYuI+fs5A8vRRY/25aCIQw2IGGYnthU2snIRB//NDRYr4chtP69k8qAR
9qE0E+cBkmS7+8KXpJKhW6Iapzx6iO6oa9rOcp/fJpIcQZIOHWy65R2Qvm6COntw99C9wZhRvX5Z
PYnAadvlQHxZ85Set7WUoN3YsUSGfXPRXyMLxD+hwSUXLpYPiaKgu7sl62fac8QmAKY7ZUyidUZF
+jgtpu6ofSQVP+5XVIQ2A1v6EBqzQGga3r2JXuHeZk6E3VUTakNwPWuZs0FZeRBVv+R68aPT9q22
fF53UUeILxxerBi3N6G2U4xvb7ymr5gtt7UR2zGYWgcdfTl1nVB32yvfE1vXm57eVXtcMkpBCLfq
kOpVj018HyMxEjNPTNbm7Boz7FIWWbAlrvabFanUZh6VZRyXg0xo/U+n3hijW4Duru5QiCmiQRL2
+eTsslZ2tjlNPd5ezu8O0VhyoZOjlG7JZUPs+d+mNvjyMl9mpRHY4l5icwCoN9UPfd0mYclkIbs+
Arb8V6ssIiwuouwb/iCqfuf8CRIT53iCB6jWoFu8E9+lLi5vtrYrND9aaZzsGCDAQDnRSAPIf4hA
K4ntJk2+0ZGAOgJUkSrKfPXFnENwiFjGBM3xawWI5KGTQDA+6Yy84CXJD8KO5EbPUDYJbP1jrKKx
WmAW1NwGbv9N4FP414PMKCCdM1seWZO9UzDh12d5lxLhQgDeFI+J3+lOhxznn9iNyu2mRprKnRVf
j3O653O/3NVWQiLY9socVa5pILPx/xZQI27+aiLnaQPkKiX7CM+DOSevlw5kV7L3VIlnz1/Z56u4
nejdckd0TrTHICzge/ai9yBS1EcoN6TAkG3dc3yWwIhS4Tk5mAqvpiNiu7RtPK4IT/TpfoWBdgCb
hbWe26trPDXutJeRWPc/lJxoDuR/0A7+me9klwrUoTNJwOB8dO4NqCavAb6cuywq/yO4flO23YRo
FetpcGYHb+2uaRPA5Vuw9AYslzPLJrTnJCJHs6IfSb+cJWX/9jBWQFMoeigpyKto2uP+qsyadTMv
sibETG1t09VDU9e8p1115uMZesRB7pHOrEmBbrITRmwu3VJ8N3ASTpXATYCKGRfGrjyy8a/oE+S4
MH2KF+/j0JiSrB63W5O2sNV4SbT6U8h1gNAJ8VqITkW1cy7n4cPf207VrPAYqFmOIB2iJTe82zKY
w2h37xNFXP66XQ9HqqkohcKI0kBd69LgVZk5cuVm/cai0L3dXrLdH1hyipXRXQ9l6OxAieRUr7kd
gs5HME5WcWFbceQJbgRN6Bk/TPYswy0fwUdFsQRIYp4zXaVl1Gv6eaM7xoi49ndP4cWcQqQJEQN2
XPBEidrgwP6KkMxCosDR9xmo43TMCnkZVD7UT5JGMKAY1ohSA41BEbJqFeOQ17ZMq3Jcj54RUr1L
uOCGiEtOhmj2dz08c+YFG4c6tAVlyv85HyCDXMrPSXqiHaNSzhf79FPkHzGoGgG/Tai7oT5Q0hnj
woAeT1TzuWtERtmUzM4+ryEWVQm0XTcKFbZWAdT6G9yKJGjNT+fjiBZhBsSxjUolUTt6vdXNUak3
4+COjMu022kxEYAQgAX69ClwAAfDbJZihElYkEENgofT2nxzJ8xXucN5tUKtnLrXcD2+967dWj0C
zXeHZW7mV/HemOUKCCifQA9insLe/SKTG5de6dMF6+iP5W6WZm7PSlzfgmCZiSN9jESUfWI5+FBu
Yg8k9Lzcj1VmqN8xJmbOJi5MP3p2qIG0AE/MR7Q2/6yc3XbCzoEFCBJ78JbT7kGAh0vg1zzU2Qtu
xguhlXE4W3MdXa4tFgfj3PiUt6/PNA28/R6AJCLaryWjALuxDFGdsn76PYkaKvsjHt2kq6dKkyyX
0HD30gf8vNkMNc2lJe8EyTjreVIgL0UXl6O9DLYIRWyfXSuC1rM1NtD7rUWp0BQddzutvqKWajUD
1A4YNHZgV2R+7uFsYn99FEfwPfYtcpv+Q/LsDEnLg5uHtaAtdz6jNXeMfOAq1v5LN1001Yoi3aDA
SgKsADplymTMdQcl1C2ZQZQTJGGvq6TrEMOz0jeEFOq1f4kwn5mTu6sESk+1afpQlDug6YQunCbj
4cAjmvb3xeuMT0Hf2xOaTznAK1xmBmDVOhc+qEo1EkVHRKjVE7hQN5+psZIxAFrPLRimFdaox1dV
dXAo/UHOUT657+qC34HY8RvrgvlzJHprkAEbi/9YbpM5c45W9sQ/ByPC5MwMuy5uWOwesxolfnc9
LyHss13bozmkdkHWzsWtvCMuhaJ1gyy9TnhZ+SPT167Z9d2sMdizWjg1IP+680fgCZjBOZ8W4GiD
z6VMShhxVphxaZwL5zgDsi6CDFjtN1iunKGbKLxs+x/j62dIsKN8Rpswpj7bpPEUg6RG8UtY8Zsc
Kveo6SggJX4pratey/8s9zqbMKzaB4lJWcm+TkbXl4gYz1WXEuCwTPMpI8SQuxVK+KTzQkKE39RE
Bi/Bh+kXYcsE6xgJoxe3Z0hNSofZBlNIFD+/yHi/Y/CUo/8tSKWn7p2djV/KZS6XGTOOygVhrhXN
6Oowu8rfMDsjScNwoA3+CLnsmaQ7Ee8maazvKClI9rOQK7vaQ3WK2dy3RwmWLBosH9hTEszmKjG4
YtG714gSpmey183smzGm9Zm67C2AETEyh3ZAU46wOlU14xCv7Q6theuvxX6PriGU+d3q2qOFFqv4
u+oNYplPv6N97HZF+FWO01myOm3ZdE64umhXbJrqGqj+RHpTbnsF7BTa9ZrS1i27e3M5DfFjBeNL
Mdmd7nmlP8Euos5okNM2cWhScDr62S8SqaR3occrvnkIAuO0JXfy976LSSW8TO6v4b7rUb/L9qXL
hjx4Aw9uki/2zZ55Iz1SmMTjg8V4+78IN8d/ZKd2KE+bKDaCaEHxEymiD3aW6XX4qq1rPpxADSic
np8dY+jU10Ke+H7pf6Xho0Km0DgC7irqYjNL5q+BoVXoMDlGV7V9RVnoxcHqXDvPBm0Liko98Ar+
V+OFXw230r6PRV/Z9avcmfctVg0wYy9FhGAJ7x6n/lFo81MlNIBk0RXjqB5WU9m9+4hu0z6kRErM
tIsWSrLmuBKOTd7pL/xuWt0WFx+kbRswI8IPoDWU//n5FxphACxb5125VoR7QqycJ0GBpn3xO6Zc
q2sjXaHGnxx/j9hQQj6pf+krsloRnh1HBEVUksdAlOEWRrAiDP1wVadRwt4empdMw7m4RQ/xaVi8
LmGQC2cK/s8LXwYmgSxrTD91fcuHgTnSnIZXGTxTvsO6wHnpAcoIpDfvqymAMpPaMig/+F2a7w3I
xT8dLbSN685lhcITaQjf9zqm+Uhn9wbxRpBU1kvQnkDOE2rs+0tuf0VJkC92tMAlLUdX8GUAr2Vl
ZwajORSAnOlmJiSbcqrWNgCxZkzMvAdINGcGvUejMDtNLERLClgtk8c0wU1x8Uh4KjAjKZPIwWWr
pdoy8sWxwML3E+NpDsFeOVCMPajZJAmmadjbU+xIKYv7hqzkpdQu8OS7M6MqCG27B5MlB7PH6WgG
DVxzcx+jcHhcW8e+3hpFTgWoLL/w9EP0LaHWjVXKte7PAid6dSAjbhGoe4xU9Wsx27AzHAi4sZcK
qvsSGzPFYQhXWrKYsRPtIji9QiOA2hD7n8jiUB9mdwT9iRjBV0Cm1AiyESmEv6eHciUg7Nit+lX2
iXE+70E1ljz0RJHr/WW2rm88tnCIaJcR995cTHDvmGgfhUhMW4ZD0AHSM3o+K/xs2lt0X1Zt18wM
2LQGeusxC7B2R+YRvLPnEHKJzrjZQlgITWkNpoDgR3QOFD9WpLBzWOVRR0bUi8R6BGVJ1u33wsTx
zVsxvhJ/0u3haMVNn19ZbkcIK9rMJKl5OVS3gIMQ9Ss4Zx9sgp5gpsduC0Z3Eu/4cRetMgyVKJAS
Y8vVRYIdQdShZO3yDgSgEnmNlMeVQUgc/K8KDCPi+IKLuUJcfCPMmgoQ1y9DLj74U74/sIWuhWsJ
wjYAHrgLfnKWB9kGYDJCYFamAlGrP2K59wo4nrrdxBOSFRucXeurvldWqmo0aQlmDTHZGBB64Wxk
SepHtH1FJfHhViXY/XUOgQ8m6+N8u3SEsJblZfA/aqkQTbhn3/f2ROACG6FkCnLv2D3QHJ+GTe94
BL8Lth67O/fassCH+yUwOCcc9tTpPEgXVHIcWSRg4li11r6HU8CLnOQbhxoc9hq07ePmYO4Uh2Go
nq1128/fUCkDYOMsPpTxSGZgB+xoMi3PwPlZPA2Bb2a8p6Xi2d7CLZGwnoX1xwJ5i9KodwFUuR2k
0NMxYLOQ7488Afc6SZOJ+Vj+xumnDg9RYX7gyEq0FAovDAUtPDXYcwHFk3bp8CbSl8K3bme4lQwj
BKPd9ehdaQx5Ph6yxKukSZW0pUW6Zq1rQnowR4fgJmuODPW9xHTAHg53rz4lOMnRa7P+ah2l90zS
dOUGUZVGnKv816rN7qjbAtl5PK8bfjzWaI063Oo2nl7e2tOtD50SqG5adr8xQNBWBm8p1Cq5fH5r
EJo0e/xnYLdEmxJ5dApCY2xmTZSMXtgOsrjclyKzL51kdAthVYiufa6VXiD8/ntjMa/cEXR12N71
Rw+AjExgaxIRf7nq8rRziBSrOQSQLytbhdgLvfYqC/B8WV817vR+299gdlHjCexZaArVlRawq0yp
yNjCe1rA0IFBobF85K9w4zEGUoyIPB1pvR/BS9WN+ZuI75Eg1GCa8AvGwe6WHTXqKS4FMah/FpBo
4s52r3fjNWgrGG20erWc1H0D8xTHknddqei+bbDhhYmCnACKCcfKKP1pzzAQuYTV3lYpJmFA7IIZ
W4ZALXO8bEk1nXKlw1AKTVclThMue0W5ylKFJp3OTGNKsSU4HuxHAqRaHDneCao2AxeGn2nHe/SK
je3oDVn7Hc39wJZbP1cpF9pXCVynkzghQ5424cHUOxtXfmp1Qf3ocIPM0qE0WTNnnE6utqUfAjEv
VHtvAFR/BuwAb+QsZx8N4xx4PkdBAKXsJWHkpYb6IlH4VweC6aficpTBTr75oRdrwwf+9QAVR7hf
Mh8+rcrqdFuiw1MmsUSDkK7CcGW07RlGvmzkH1ilEv0fLggNd+5xsvWQsCC/gIOWkTd1/s+nm2EZ
V5TbrQHyOXHozPfL+sX+NtK+NJY7u0ZBXdmpGl7wMWgqY8pMTG/W249Jj0QZjS2StCFYLRvfLPQV
+6XdzlVI8YwH3QJURhx6SVAfTS9M10qEat90+G6X/cStdHhbeqlxUiBztJsT1vQpY7EJ/GyTwsxd
ooXbZMFgxt60EiHIO3ZNY6uCKyZ/pyZZ1aFHt2Q3b3syXZ2cg/I62tS56Lht8JMk6fLyVlKmMhA0
fWLxOP6d6Ys9O4Yq9U0UKN2WvtKBAK2qkdYK4Jm5DDIFzcqKbP9mCXLXT1OWEjbV5gsSsvYCWkAH
Uzox+E/zV5Di5m4BCtSMLGVzh93g4OXWaKHOmWtdWNOgSjYYLtE0uTJncY0r2Bp562FgIy2nqh3T
WSMwemUwbR/w9DIIz+8Racu92OB3CJY4UjUy/FP5QyeDudk7vWsYek69kLfs23+lEBnKMs7tbTgF
OhE+Wa7eN/WO+CiXYD+l5RzAdqiyPaAjojUXI8oEoopCme4R7CRzjrMxNjQ/lJBne9ySO6ZGSusb
PZ4F1oJXdh9ao+4ZsMo+uq8N8M8ntKbMipQQ6P/ZoKUeohoA6g3O91COOmiqr68Tgpc9TQgkDs9x
taeAMc1wMlxKDD6zkFceopYXO/ywA4nhahV7bhRh7cvCYrNE2tq7r5+YgGLusIPMBcIWuJOUwBea
qoPy2WXnkr/PJrHuPF4f8ZI4eHL04cEN1CIcAHncDWaV8NYjdPhhjdIDAVnSPfpAitiH5NhRXDt2
RRJXgUAzR03zWEoon09N1AiSSZXwaEB9C/UX4i32NhLpMPhPa/ekCmyukD9H822gqWms0wNsrJOR
uY3YDsLhBAm7bEDayj8sMvv6/Ufd/US0mk2du8q2r22Pm2aLYXXYfFx+s59udRZ7QKQlroZYOjYX
y9DtoOPmgSl02LXRl7MBLlQ3iVWgdBQX/hy0ejfYcu58L3PGlaM61TfMzXo61ulP8wr7MpAJe0Ut
8uroApBg7wotIsyod8ZWG327TBr3St2dKTV45niqmDWTbtPBw+MK5RcFCYZ63hpbRqRG1XSrUtcD
xXyAF1kO2FdgRUxZ29mMhfwRTYJFmkZt7m6VQWgJ3mG9aVtbsaqT7wkqcwSIlshJH4ILPg/vKXj1
yVLIl9r/bxJdiX8T1JABIFB11bjcovStL9vrrmMgB8TB4NhNCgc3ggpJYyeTZzpIhMBhgsrTiHRy
lPa3nwZV8mBXHe/Jahf0xZ5NYHDUaeUMzyGiSQ1tmDbcJ+zB7Y1rByNNfiLyoxL0B1yCoL5rlwKb
VRnuaE+IxN1VVeDyEkv6IKQcYBVNu+yqdxUx+Edv/9ExiYzTA0pYhf9F2mmuEPJ9C1tk/SfYrdCc
NI0hm4nF6KUqlNdt6N+y11XHblbFqdkd2y+JyLRPvMsRIvEYrbNBuJI7AUtw4A7kkETAHcZwQ129
Sa3HbLTIOK4uro4/9foR1hwmc+SYaPDhKCf0rK4SKRJE5KPdIcHGeOUy/YCFsz8wqfUYzzO8xMGU
NMq0SahvWv/VcIWTzaXbk03URIGomDD5cWKJLUfPnBGOeaoPcegknsTXuFtPi1QsFQKZnPLPRHS2
O0Wc+K0Fx9PIo4hbNGhktyyjYzvykfyJ4XcQxwtos3l0izqeFBDqpL9G2IAomjUYaqgIE5L6B/lM
Q9SoaqfSvilD8GwrGUgYpkFjTtGuYaHkNZw0SXRl6nJOm5llWX5Pyhilbk0h7PLPX294dOxTqJsB
+QaAcvL59LikFWDNr0Y5ecSVSFVokyBYeNPqU/jydMDN5NWfdX4xQvgqJdB+3ytYnpO2/nnV0tsx
k5/jZJqznkcPGdGYII3jNtcyDioPh3Lwo+Uwg21ZxZbLiOZ/6p4NxbdqeOR9PNWqNO7ffFsV+wAH
KCn5+phKbsXgTLvsxipqJIahXDeOUbbBPdx4Pk7a0wksPFro91RgWjYSVqVwH+gLoOP4kuUlld+C
FFzs1oMcBUwH3eSK6IAt2HabAeqbDFbX+jRWzzocSc8oKBwrJ0G8hMj3ICHVStRqzZ+r6qmuuyoA
eDjZr/xcfizhdFHU+iltv8bTk3mlkk9E+j/ONRGUdlsqrD//cMSBrmKcODPUwPWyVz/TjPoaHoJR
kFRS6EbvodmGm9XhDoxy4aY5oxuDrSa0US1meltcd5FgAFBPfkhjetFteBm/1L/HsDSIvwJE+81l
kM2w/P/1JvMrLtR16o4Ct6Qf/dIKNpz9KM8hcbCz8eMn9B+9MZJPgN5lQQxgSCvqaTRVgN4yc2wa
C+YtxIsNVqnOLF8H82xxmvR3fdLd6rfga7MG/YIbkyQE7nyJ/FOczbJ7+iVhweAn/n/pnx2TQ5eg
/PMWuJl6+g7GCh2mH1raui/89m28wF1s8rglM4GzHGrZZU1Oc0UmyVO3Yqt0zLd/2NYAmGLMFDBl
PuDTWR/m5YAVQGtBhIFkuqpQlp2qA5LVtvGdhREVCtbU3Arb+8ccLyZF0ixxjS9o4wnyob4vxgAw
IiEfk06oJaORizqliCmI7p+QTJPZRFZzh9AwR8E59KHaGE9J+1Cw9CwLoumCRHFhWxc81J5pGIka
kpBZAkBYBSdEGM1Jht6JzZFcHk7I8aKjc0k1UWmIPVARzTZd5/P+RLmEH9WruUhCc2iX59pw0iB0
ORVhsJmN8O3hOssWG+bZt3tup+DVDbXDQnj8tWCyPFX2Z2Gcs8d/MnQ0+IHnvVP3h5NRDXMCoXFB
irqUYhoX1iVcgdkfjTH7Jp1NC7oISnsXzFGbHcWgtNGZ3kv12ZG85ckpoVHZ3ByWN3ynmvJGALSH
PoGBCaW6hOlPO0PYWA3q3xW9oHQ7/Zy0aDs9Kq1ndQCfa3sPEpQkKoBFTha/1/z2T5GhVTootuel
Ht0oYLkRF3T3MbN79sZwbCgXdcKF845BmVFxMtC4sFVYpUjFaJmf3SsAU1YyaL/nanJ9JYvSRZin
zv/AFu72796CO61TPjBtG6l7YX7X36UP08VhU9/NHXPUzkIF2kmKZP3/H32Si1bUTgqImvubndmQ
AE1mCWEjHoY4/ZS7rXbMnwfIXF5KV1RmcsqDSq7D9hcjZpWxwG+z6Odwo7uisriqh0kFyDNAXq+a
6+y7rEgmyYu1MzYhxDSRafugDxJddnyVu4xVJSGKdfSpU3vEX8oRT9SnlD3q/vdr24LVXB+w0fey
R95saNC+BnT3NvL1N5dInVbJ4WeHgD/0tAAvoyr/hDDiHbQ/UtPUXVPebhQAZCxPN07lBAV3CxwR
RAftrjTs93uQBoqoIaCSXWkD0aQ2Ze/0tb17O62R26GSd0k2SwNB+rW+pZaY6ZuqNlfpIyq3B0cF
pBwHtsG3xpcBXo1AEx4fuuGsu48ZmCeDN7w2c+952ZfeVtQ0ZqthoKqIw0vGiDzSk2fe3+5cjOs2
rS5U5IjzTx0JJcOuqOsOR5AGIrKTLal/YQ4wbU0OG/6M/iOVGwyKV8XVYcrKzja6OceJ4rq4zAj3
N72IwwXFlYcEmApQwUIso1M=
`pragma protect end_protected
