-- (C) 2001-2016 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
Pj2bVzsy0CApSTbuh0AMN6ZVE55hGJ5rmahrjTHJaro5rfrmz5O8WADKrT9giLL+IeOFw6GADipc
bbcDJfb6SWoRig+xNaK1Lp9YDawIT5OTUzvL0Vkupfp887pIKHENn+NwvLjhHp/oIRyz1Dvig0q4
HJa+BXhQ6AU2QgjnnNQGny8SICKE1xxjtTAFJ2l1FNnaxFaJLSKfP9Rh8mLhg/kG+0b0E0BjR0hY
vHnEsQRA0LBYpj97mxmnGElOoyWiy0mEgkI9/ZvB4O6dhgj+G4qfnVuLvJ1hykRBvHkhNW48ZkbE
zj+LullAZXAf5hGZds7AY7RHCF81byuEVV59Gg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 4848)
`protect data_block
P0FJ0NqHZoyvlG904A2lE5E7ftiSQP6eaOh7pw5FSdc1qKyMjj/jqL9kmhRid3MTspw7f2FuUtYV
wwG6aDnY6hu7uNbqhSu/okvFOmXWGrJj6byh8QHpoajJPEeQvmo1VNxie5fq+mEntGPp/9QH+gHp
XHYOk1a3NI+14t/BOEttXWNAv+Jtg7mYuEZjljuny88we4lCw5fqLfU5YuTmP232itiWMGCIeU2l
v5i5lDr3xOotbt9ojpAIn2chlXTQk0UA3AZxCkGiG4QuhZYlJ99+PglJBrcnnETSqnOC1XB8rUlo
yS9zBsCVZPV6/j8EOcI0QqBfgGnd1eEQ3bjLAiGDizMu5NFH5FfBb8y1j2Gv/w1vD8eN7YhWt5Ma
j4SY+XrFcWYZjOkbwsLIHScxnr2HxPelb67r/iOhYT7zYfGOYrnQ77yP4xuqRYou0G7VXklHy8pi
MBtpf3nL5pBgvp43kVM5WiKGafQ+HubFfZVsPdR35gTNPJCqSxZVPZKfarK9QQIyROO59r/GN6a8
YUn9/9SrBZsZVyIRqDXp3PEdG7jUxWZJ3AbCQN4ZJdT8pEPRmKs2RE8SFuc3V4booxOVFmNOe1jq
ITF3q3AgV//IhARx+f3ZHNDJAP36II6miaXuny0UFL/lCmT0PfyD2eZPX8t965BugSeDiLCeXIHP
HZLkMQsNwJbtAv9yk+q5rNWrtbq5ZdYynrWDydUzUSk9hTH4sSYx1jvQjmtFoAdgfXC77rLvsj30
qiGSfpcDzNKKjlqHPcE0hTo6+R8LS8M28TvPtYdzlUjcwCOAlWXrPkNs9wvkFdDjJ8jN8rcOOUrx
Ek++xtWNoIBE51H5mWbRMnwiPTQuTzmNQJ0VgyH4Rhu7GE8609qJ0iiBn/gv8i4Z1jFCCAPekC0H
QJ5nDQsfqt0PqGjr35M6J4qdQDUPKylCMQpRngMsgPh4uGpw6XwUoE2GN3ZREWDNNYkzdn7EZOMZ
B74vHdHB1mmJKS+RnDCsPdc8T4K8pCiVfGaNuQPclCgw+z3mjXmlxjJckVydGI245uMy+f9p6GXA
jCtV5/3lxzx/50LkpKO519M3O48MMXkpScJs4iOBSjEkC5OgaILom/RF35oXDbi74gQpv50tF6LK
5vMpGtPGCA6MJ1fEQmI8mmB59ryqDCPV0RCklj0n/fYBzg/wWT1RfBkzwLeolFxWbl55QP+dHecv
M8P4CTkI56S+lwDUIp4GMFoxWTE2Z2dudNZF87q0uK1iGRuy1djRr6JppcjuPUmMwKmpKdmyfTRf
IpumOEES2v1/5zjsR+yprmphBV6IEdim9fXpYu7NQyRwPr1zp5eCgoZRrfrctktDMUkHvdf5OGem
mBH8R4sUFGoGRW5m1Bf54g2vBv22wtZvDuXGlpoleD08z8NDaHWe3CrRNJNiP42uLZI5rkS1Pr+R
GksYnDQb6cLdct7C/sMpxFtveH26WlinLTKc+LfVcO0iYvvIcYBaZ6qwQ7P8HefJlC48OBud8XkB
R2vXol+kDRO2PyYUBp48fi7QR9T+nPovu6NY2XlCjkezvOBreQXKI205cyMY9w33RhpNNpl8H+TB
PgqQnzaFu763pwq7DWxI2CSEUbwSLDp8CTaDLuHAwJj10B8/TaUOxHWwn1/tRbp96PeBdXM+0TDC
KBsvvGsEneb3XmyNOAev0ZsmEYCfF8XlcFMTBj49UgbIqblq63BM28YpxENJe2FbYCfsDSNWbP4L
2w0v38WJQJb19hmL096n7QDfJy1XoNQnRPyQ0vYW5Vap+RNn0Z7QSdPVP47uS2bb/XtfwY5wSW+z
nnPzs851MgUfkNWTatt6ifJn9GVh0gk3GWRUfyrc6c8mWDnh2zXrG7nU5zOsoRi0/EaNaDmYJD4m
MeQrUblDtQMcemv6xfGrE43vYNYPuyTrblvdP3yQJ+iyIrpSxkX9+EAfo6PwsECYO4xbjUPQngq3
TwsIftJiX+y5AsAe73BnW9Y7FdFhl/L07yYXT+x5LCiM3xCYI8ubKblRhrvGjJWm7zxzBUrwK5m4
EP8f95IhzH0fsu8GG8CfMpn+yRN1yZBGCajUhZWI5NdPUDi8lIqnYYtl6yxeh4U/uyQB3nKuA/6L
dGG798D/H0xBc6cHhxB+I7pHS0NY5bP2h+BzQcWwI/K5U2eIqzfKFLAH6yutQbwDc6AtFwIMRdzy
/ktVwTov/Aow13HrvXoUvYmZTxnJ5L6QjpKcw0zVjrXyOXce9iy4X7rgq4Y9jebI0A7B7QTk8om1
ZMNl3JQ293DTFgj8Dbl1GgAsZScUifRA47tHkDgCX0Tr+j4o2mGGX+VCwY7bIhpjQqe4Sm4ohciW
QfqGLjUsWjhSV/PZTsSGZBVnh8VNs+/Z480gvo9QH6xunSCeLlcjsr3VIgz58rc4dPbpbPdxBUF4
QL8ui67M2Qk0ZbVodG/h7/zktC2J6kQjhIY3tBQfr6+zyHnR4Xlzh6UFI1rffuzPfinpmxuCHz9b
OutXoROKN6nnlyQlzcAlFtfG4dVtio0zU9oAfxXjoSL1NjxTqErA046rTZSozT4PzWluwC/+K2F8
M+CajjZxsDlrFGnHPR8Zt/8ddVv4asziVcpWY70AlI90YkRUVb6rlW+NJg+MAJkjm6dZPJsEtA7Q
pElJDPndtoRGhw7F8NO8Y2RLvBRc+wMjAtwZgsnd4kdzZwrF4QdwLm+ZVcxnpQIe8KiM7XD2YEeS
DXQR5MMdGibj008SGVgQxpamygqiC/cNT18OTrYBXbmzYjkrKszZJdXyFJFnUTIesy8z4TQhGZBS
4wfvQU+psIu6r/YN01+ogvfsn+e0HWnB3+VjovZb9cNETYjdYFEDJxf769VeOvAChuepP6KxRLKF
VijY2BvKr4osE6JCBoOjFAckKoyPP8MoW4RbcV1KR5PdZV4Jpbu1aDZVKsFR0b/CLmQBxjiYbs7K
tD4kK/mbTiKKGVhjRr4+ZVS/OCLzCQpmBeJMW+bzk3l26Jzu7RO9NJjBScPW3o2bd9bkYsMQeSqt
s8ENTTAF76L7xzGlTSpB394HP5M0IO54U7ujc4qu9LQSfMQjjt90YuCpmNAz+I6N52zkWA0G8nP0
H6nmOv4Oh/XCWgvUkFjwOnbdVRIj+8gVw7+oUmY2qdLnihCQnUXJGnP+hXfjR88Ck2mZL4t2huB7
TMLj9FtcvQmwk4+a/056BtNxo0EincLbNzIdqzRv9qMFBiyutASobKDTaZA7+kRkk7DAH2g6dDbh
aVPhfNsKPikf4Ffp/96RXWyt7weHK5j1nwTGnmkrGUQ7nx4PVULUEDNYNwbGPd7CF2XbsqlwBqPX
q+Q5n7huzpHi341wepFFJlGG+KfO/PZ8TCb5etXH+1iIjRLTZPXGJIVifjvrNuWCLcSWF6zkOz1c
cVDVO4K6Y3+3EfBp6OlKkWGYDe+3cMLbUAcL8K5KWNhhKDww+z0OxTSJ8KcEzdTaEff52Dh/7vq3
4jIxTGcUP4+ns0//3cFNp4zuxLBqYOg8wo8yif5+wWtkUz1vJAL/CdCssvV+o/65E7z/l6fgBIXs
r6Lr6idjxwvdpwUDVPVoZpi3gwy8Jij2Qi2hSEQML2o/k0vDpL900iewezae7jmc1trp3vyvLxtL
MtI1A0i/9n1uChCao1T98sji27JLtfW2N1w+JXoawcyuFj+uoTpYmnZIkf0FL6PJOcwltIz7/fO8
74yDbzQbhfrHn6bt5LerfiyFj0NMdOVWwOQ1ul93ZZUH5N20zclr6qLt61RvIBcEvKifk0OlE4bL
AB55NWbHGzRPu2UCZg+qGMgaapvi6tHe1n2Sz9w7NIfYUBRG9EqOq236OSyBCtNkIvfEcPRKtx0h
K7nIlvAC3phv/g/jnaXoEncJ4YBqgjju6zDUuYa7tFEeC95dNx9hlllq6pHnPoto50SIPaz49pBa
xz0gMGUKJHxJ9aHXRBuUeXOH7jJdvMMq1ljGHcC3C/lSFNooFaVZUVYThzE/+4c7mfnmPr3viYkq
Wt8OTEOdFwTJs7bY4Y+fDTDcHhIPa4Pz1Ut/PRBvM4KYgPj+DxYkcUOPH98y1QJMr+pKuYeGbbBm
3rMWQmGWVjsKfASNtbwnOXH37uPuOMJUZn0sQCG1BbSXHQY7dMpLTtxV4Tylbq6nNds5rmt7B3U4
TqD2YpUZlEqk6enMlVRDvBrpKy+FHKreNxv3ZAb3LMW4J0CtySEOJJQzS4Add+ZemGTt6TxxtgXC
IPtnqspJhNsjIhE1+hF+qGgEtPsRFbkeprWxv7/gdFxl9oVYlcC1CAwILZ22pfImsC6L1Z4aZ3jh
iFqJetl7/EP/k9crS8f8fATjK6yx0BkiL4/3WC61lxFbBFqCYrnOXgvttFr7Ma301RY0sLzNg/9A
AaHtgckFqLYokrbmCVw1tzIzVGcQodWgh16p/db9GXmBtD6+PDEmWwfHdtMCK/Ck+XPmFbF7JaNc
m29uP2SjYwnMq2GQI/WjA5nsnGsoR7cipGlm88WCOUvMSwfhJ6CQ6B/FboZ+Trzj2SVZ6m27S4uV
+rdGL8AgvxMAKbBKsErT20FSoxC/4siH7aw5/NdRSFWeqFPijQcvrdssFUurVaj4Jhwoj949BEea
l1EvhciJhSwj/Mnif4JtAIqHK4ZPZRTGS/JUVR+eHNMw4yenaFOkF7E9dgnmwnT1ToQnZwBOJYvL
oRxKmcbekWEyvsFp6UvO77535QKxR0s2RF6Pfkt7NmyU5gtRTdRuOqAEIC5uZTcZMGCsDC3b4el2
yWEmCXRrOBg+/BavoDwxhZq53b+VyUiCgAgW88sJlzPAyJNFXssFbDFuyqlTNf0UK6hqrfhIGnqx
18sDz7hMJZhrIkNJuN/i6bWxQJXVJRMhLCo8QOsdWSli/cbotkdzKHEqWPaI+yp3g4Fv569f1vtC
IE5K5VZeBLyImgZoK4h7rU4jPMn8uuUeJjWfpx89RiDKsfOkeAq32jM9OdOLfZc9qio4ZbWdlwlz
91soKo8E3LVbUcyYd2Pk0EAOJ3BnKr+EdMzzfoyF1liQA1PA0L/i07pNU3f7X3t3DhjqCIwvUmqX
SzRc5tDba+byzuPoPKo2+mlJfNhC4X+2gPE/PDkb8XWwRV39xq5uo0cLlKL4bT0M8e0d/EoA75sL
rBX2zN20+KEnjgKfMBImaKqE7LMiNLdhZYm1znNBQ1iH7MSP19FX2ijQptnXkNTKqx1lRCfrJuJR
DY4GtjF2J9BfNRGyJl85QqZ+gAL8KdcbIKT8jmGKnv3fG6X/2yPryiKwwmAkg3TUk6GlgZrxTIiJ
qLQxVp8BfReehGbOCSlNTHqU0FoM1velOFApY1tzTb7iiyN+zoCn0fUFxgpJvuaCI/McXhvfq6R0
dAuj1fDlG3cAyPDxf2WICSjxo+/RaK2eX0UXAeTfCoHLccEWp8dT6LBMk6NfPilW/h6P6jg3Los7
H+qQGcX/262cfC07JSujKDnoWQIl4nfL5Z/ApmS5NPdzrFZva5tbOYCbQ+hGrcoE8K1Re7ekIHCZ
UGAI54I6Z3uBZR5vc49UkIRE98fV4d0hZ3auyR9tuEDUMdIBXll96OOITO2lOEtx6sEv9XQ2awrH
CYgXzkbDRukwbL7VKKNvLgmDBqZimcVERs65QYLcf+30ODLWIEf2G6sV1B0uHL0hqaD5bSEfUVh5
Y9I3rfI22jBn0g91D0LxiALl/YIIDiI753c3fZDpQKx9eC5gLpTWVJQtR4IxlzL6+/NLAGPOi3YV
SJ80A24FYUMGcL/g16IRIvD3zhbDZXFPWzX+75aHheq4LU95pX6RTSUqu4aNzmXc1FEFJlGTMXQs
TFd3b1pZPJ9hvN/XF7lOIH/XWI6WqWtwfPC7NdRHFgJIAP/gLq1lWRwCOJfLekoDlRLo21PTArnO
CEZM3xkh9fR7NME10s46oaGZyUi4JlIvygcs3VFI2ZC8s/w9K9VShb2wCPaSu28xU2JClfXkUwa8
MNurI3hC8OPWqW+1yLIml5LnCMH401WAV8kRg0RSNmFyfFTsU+zq6psME3wmYBDWeEb4bsdbq/s5
SQ7HyhTbkz8ring5yFZfftZuU6fH5mHq0E8fawT/X7nJF4roYzi8HjGXID/yYnR6+GgKuA5+1jz8
RLUW1fCcLkCjW4FQ290v/GgFM0oOUxVfdCGohjuXBCHZYuyycJF2dzncbdQ7wChEI/zUMGHE/tXc
9rJZfW36bRva2Op6QwWXJBq5ieyCYFlvUlCyt/F29bfDE14oogS+wALARYGn1glG8rUagD+8IKlf
/bw0p+qKHc+xYjOzZw+dtYUPMvXD/Wf5RUAJOTGyTpQ1B0awjS5B8a3pggWTHvtS7z9XsTCMCIP5
jervJYwXeAdyPH/cpQhhJ3QTJm1hIaIi2Nl8sO8cEcYuIuOxptaBrM5JpHqgB+U5wBDqw07AlsGr
dTNW
`protect end_protected
