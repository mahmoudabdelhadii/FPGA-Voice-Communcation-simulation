-- (C) 2001-2016 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
lHgBxa4rBkwepDjLQcOEpopkNpXuimKZZZrqaobyeE331z46YBwGQcujJXSlaWaGLtfJqQX99CLo
zAKrRk44XXkVHWH6w29iOq+UTl88ROY484ofy2JBO33AES7gGI5xEp6mRGN66hKYafp9O96xEj2l
5lu5nrBmtGIZ7cElIpB5ntTEX7ELubsaQGCz0Rqp0gM7tVuVPCj3nua8xs5z7sS1Nr45hrAcy7bU
ROzkVGNZ79uoLFLZzc/pHB6VE49FePxzOy2OB0fwJnooGdOIhdzKdGiqp9VUcUNNS1n5G/Xd1X18
CeJHbN3mbS48xefrKDPoFk+NYNu1+jnqIeNilA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 13456)
`protect data_block
ghOqMTy9hGi80CCpau6mY0t2JTyN8TXBUuTNGYgMjpK00xL36dlsPeUjQOOEnUvV6JPNHfUDt4gT
B3QoK0TZHMKjoUg2JFLIC9OBXFJs1iNNvrJRqx4OVov1qikCGdmSFtMWK5gc699mXrnb53VMtJW3
fpQvpBXR+YEeAqQ3dMxn4PQLPxYdI2WVBsGDH6d0WjZNbMnLrDk0OFjdymKtj2lP07GGZx8GO4Zm
xPn5GjYNHEzf8d+BaE7aIYFoGBg+n/b02YXwlG0CMiW6njzep+BKh4X8KLFZgFKxQL3OwSZb7B0x
zcASxVKR3IJMclczmLR+jTw8rFj45XrdsdLnMNGtjbq5Zyok5eiMRmHpKcVtPp7bPsiCysjM2/vS
+wNKDkYW3OuZUI38DqWcN0AbqLNAxaW/XkbN5WfPN62ZVAb1GK21ATLFh3EcPzppP7pl5uZQFUJ1
yBENIK03FGBz7npPJuSwmOquDWICgoMwkBNk/0kZzBTQbqAPzdAQJOEwoPr05q2WGXYwrrbvB2HK
SMmbnvo9+RPfesMM1WdmdYogICtR7L2/HfQ+eMi3FyCcjOvulOUJMAOpPdSxCmfF2Qxc966UoC7K
OCcLK+Pyw45BtuwhXGgeVClMfz3GD8VdSavhIzw9pe1J+0Xttik9W1vbAXodo8yb8OG/CWAEaApT
iyX585QRCnnaT+JTO6nKpjchgRLcg1MuTrMMAJTucsOoG4uMjQpAMTV/5y1rnxbOV9mTgEX2Btp8
ANeS4p71lF+50aKk79LjGP/NRHNggmcYXlfYD1IRwsb/UruE7uA7nI4K/D9e5szI8tG7w2iS/uAO
rQaHMySKyuhci5I3fZ7vHnFh31YRVoLeCIp9ikjglm8pHYU7ZcC96i85MrTaNYb+/fYBh73fhnCo
UO1FvPd3AJohWwvU7ZpoKySm5DS3Y2nKCEzkEk4SDLe2wlgbwAEGbot4cEwfc7+i/m+DgB+9hvFi
Hr6Z3sf/+DYAlEV7S55HDxUCn1XZloMhu+zBD4nRLYX4tGMIL1mzEh0MrAk+t1uGsIKaZEB66uVx
hPBHYEdth9JIfSgiQZxJiFpNehxsBRuZOS3P4oOlJ4oNxwzSxJV8SNkakxKKRfUgDPNwwaB3aM1Z
1+ts/F2dxXKP5a3Iw3AGag3/q1j6yLEY+ONbhnwRDOW3Umi2uhGE9bfEINO1cWvE9K8fAlS2WXML
10vNsC/7koNuy+ovHUJSuX7vJrScDRCrild5JBdqrY0X/3L/sI5Jac5f3siPqgy+nESzLwg/+hqV
lxFJc/+XRQc1p5kS7ILgQt/ofTBnCvwJDVNYn3MUw89ibYQc8ppUsUqUVO4JBfsddXE7Zay8WNTR
l0KPtvEYPXsbGeTg4bFxthjBxDGzdSFN4d6/kaEirMRzznSdGUh5UN7Xis167zhm6FItGAIbHFW5
xXpbOK4r6uS2pbwD7Bi3UiXxsPedqcPFFlDcnNKLjGv6XvkfwGk+uF6UqTSUrRkG23phhRyBo4M2
J/9L73fK3CEacoBh/nandiLfb/4IlvnSPnGSmN1CwD+1U2rerSkky2WeYcYF7myjKOOfTgnPRlta
O97tjdv0I8jc30gUomsqnNnEoc4nND4qYpQTjbX4malBA+2/a+huKPRlDEZixBtIfMS+oDyHZVs8
r/8r/+rO4Vl8NRSE5nO29CnPWbLq6bNf+RHO20kkHC41PXMr0hYcwOL6rxaKqu2cp9knpKF/HeQo
zn5xKh9oa90+GElu1UpF4YIcySY1gA0oistoZTdn15S1B8IHGDBMOPdymEWVxAhA2QzTa54mVJ9q
jrVCv9nurRkcgpGsDI1JroKZgZ4QyeBOOwkhCk0iT6Z9387P8sIVMV0/uvX6Slbh96+dKbX7t63C
DxDKVchI1jGWxl8cRO5iAkV/wiwZRQienRAlhtmagmHO7kHEPazE2zbAG8zYGGM47UGfdB0+9Vas
NMVbfqqLMR4Z4BeTDiA7NQioQt4W7CTaxYUSxGwO/DSCURFGMffVS4M22irMHcaAFBwlHK5ir5UD
UEGbGorIixe9S5e+OwaY4eoQhDBkQeXBtTmQhBxglmgSrgUR8U84nBN4pCpWsn/eIGJXUtNmQ+GI
Sk5LDO2ss7q0dcCEK+jIeDfLWoscUf/YB+/+8JiviXl2peX1hZF/b/yX4MRN4A/kW/AZBb1Eb+iQ
4CiJT5AquuY8aQvduJrDWoK7MFzzS8X7jHR9yRQ4NSTp+lj/shCgLFUU8pZ8Ql+X3P2eLQoLU2Q6
EjR79vGgjY6+bCmJZfdleRQY5X/GwmTkBupFtANehGRU7KcG0ZpJiYICNo/VIgnb8rIeCSbBDPPk
8hyNEMpoiSFmbfBMtLowyJm6eIHC8asov4fUW6hfwdCgjpeemCq8MzFYhGHEVJ668XaW9YKRX9w7
hgLi0F9HJpWbgCLCnospvwv+xMdm1jfGlbKlFALL8J/Te0IemsLZyk7UQnGDg2uB/mgQz/m0rmb/
bsHVcZFXuQz+6O82kupcKVBX+S92N69ME7rUh7TOLCbBRE6dp9b0Y3xJ2QWMkB/pL/CpQzoTSELX
HkvBiYlYGOSCbvdVLBpE/v6UwGcQgPImihJB3B2SuQTYWYuPDpq3HDf34IV725dJCO2sWSZVdGJM
o+OtBd2VZlksB+gU1fCOII5X7dmBBbkEm9ReFhcxRmkbo/YqknHFWP7C6nnxcWZzRIEmbKwphNHF
8bUIGQHU/sWgHUzyzLEjHP0D0u41fkMbA5yP5QzphlV1BE4snSzDl/zQ/mOoVG3ZIGPqCu1wLY2r
U859LFi8Z4KmUXhoUIjh3HCojeGeRP9UuvfzGGXUPfI8p1Kiu6dfOIjAFyk1044j8Mzl9JDVHJnQ
kUH+9gpbcg7dGSTR2N2+4YTOxIf3MXMVDgvyEzrqoDIhdEQ9Hx4DuyAg0IkUOjX5o2tjlW+gu7nx
P4ThKkMASSK8cTbA2ZKik/TScGfb2PHz90OyGcf9wlyfk/cOqFLSbxs+D13XiYjrj83BXTdKXi9E
WJjK2r9OgCjxWuIgKrHIgiBspdyM8Veld5mjIzq3oYE1qqNNxi/vOmur6HbrPo9p4R1b0HLT3H5/
jjoJBoR85iHOuu1V2CyzZrceC7Am9HANdaMrWBi95xwIsXIPCY2TMLEVzX+mxll5NVs96ypBjSja
kUxV8GI5zokCE1MGFwYZ7OG7N523ZRUfyy41NiRwUPkJJllZWKRdPlgJPXC/rwbrr4/s1Jcdzpdy
hEJvuTGPJuiFfA6+fKkUBUx9GbgxKnCubU2H2NOQu/9vAIBmTIpnS2Ycaz4KchGTj/Wn8vcOYXP1
DwS2ib7HPQX0YV4TNzmCu5VQiO61EysLqNSFk6/GD55MQP/QWpQFwHFdb5nLIEk6OynSfaSUNyxT
Qb3v4fVcHHAP0O7s8u6i7jSGK92BvSx3wM5TEfY8hmG/Fw4DdixriK+uHnVegnmfvD/6lFT3kVJ9
FxINtIRNnpxlr3W0WjVUfm8n6iM80TlQmJpcis/f95H1O6O5oX3B18P6W7kNiBi0OyAPYRryMd13
I5Rc7p0Mq3JSr0uDJXJwkyBVGZW+RTNx2HKu6YZkZJBvM6eBaCVdyreLGrReCb7vZqF2j98Gw+je
1OGyj7BBmgaXMlwiJQvjq3mHh3EzIHQjV4sJJdWcxmAjaEUaYbbnZJB6hDcYkI7S8QiM1M01Z19T
V0uPnW+GgaAsaRJ4DBBvhXyKZW4nVsipzOO0yBkjbpyAWt1G0KgCOLI7bGm9J7IBXasHLCVNpLO8
bkcqnNDy+8ahgbLvDqb12GkBGjvi9cJqVin/eDtWuuvugtFWUHF9jNl7Mc33w72rWcGw7YqKoQaa
kuH0bMbM/wAst72hSsN8jk7nFPXh2MG8m6Ms7nACtV0efMNni2/7J8FAPTazpYs9rB1tAyuE8RgH
9d9iPxXPgSZwhO2sWClCN8FmHP6hzykU4uQiig0hcwxGmJ4uDk24MmESDV6Hs6WBULCfCoumLN2i
7W/B8dRljAKHDP+yQ/aWNANwtq3PmsKN2zxty1AZYZ6y7imV8NF/u1guHpmqbGoihkJWpUAu9ucW
lhFvRqxHg/yaHyl6v7ZD7HPCRrE08A/2ifE3VX/xR4O6GO542BnWF5qCS6TYGwjsWxSxsVVZ6pj6
31GUS0SUhoV8ljgGHSDPZ5Er9YuF1BvLS458mbVpYvvETuRaHMW9fULM99JYrHejom1mJ58uwkLp
vU6bmjIQa9h+yXAmvmxW3T4hE051+rtjG8YWOba2G53fLKtJYiWg8+3HxuZF1b5OP6OGYKAtFUgc
zdKsoT0UyXiog00d4cpD+rDPOEKLYjQIeEcWwCDMws1vycdBFsY07iAdpgEDZCo7gq8cXzOF6i24
AUWP7D8KgO4FwlIru0DctngvS2wUzoA7+O2zDcAZZoXdy8RjuGeUfBGeZtEp0x/pzy+oOLzpTwO7
lUlEWZm1d6u1S1N9pv/c40DGAsvd+Re7Yp27HNYAHTatQDs4GbeIEvtLBIC8O5iU6FOVOSycY1lT
MOKFdXcQt7UYM9fbouel/LY3je+A1TMqZJMUoHKcy54LKBfQ+4owDbamtZDwWdaKepzgyLuP6OhA
dv9FDCr8eu9b8+epK+u9PIwkRDo+D4TucahA3BrmwTDyp66f5HG23pVBH8nj4reqWeZqK3ueX7NY
eMFiOiKJkihoSxfksc8Uf4hjM+1awEBWyAqGsSREBy7os8a6DBDdEAND/ih1ims6st0xUoHaE7QG
5a6Z/YDEJv88lcrfX0VXg0nB6Kkt1yDZ4RSjyHYh0GzrgLU3mOOt9MBDufIHQngNCjX60gob5xGj
gMr8YlvTaLJPnHoNSgtossl32PuZsDtcD4DAANKcLfczjDM39182BrKLD65EWHnwmBpmesx9HNOB
jJsGk2iKtxY3Wvs3qNPLKTdzvaQFgBxkC+r+EYzJ9SM/IecCs/nyz1fuUiJG8McnnP6hAKvsBUtX
QJo79641uFDuExgTKdLG5TbUzBV+oAzJIkkMrJ7VFjxTN2Bu+G+96s/WpxVgd9HKRQva/kXxrwVq
N+cyFUO8xBGqH7BoyA07TN86IKqEigDEd6fmJ7dusX5mx3qN8Nq4KcZMS9eameJDxsmDn/CsUwBj
LD9kYTSVpAEWoE1qiZpQ1IWz2RYcEU29hILWRTl1fw51glg11MvRrXd5PiZuz0Ql6JCTGLEMM1CC
gcsUGKuUWxxNmKNiFHw9c2mC2jNK+ICRpZktupJKuuBnG5ZSiytrYuMA6EAyMFlFY3o1uQR/rvri
0Cay/YU5XMv0/ejbJQ9Fzv3JkVJL+cuR72vwImfUiz92NOk+ZsUW0SaSCM4w09bWb9SOf0nPjl+F
G129n1sO86V3ujJ1NiGPBgKVKanKilvgOCPha+sOZCPjDDh4rITUSYNfA+Wu1MuQCU3w2RK5v2TU
u1yTQsJdTp7o0r3auSaOwlUwwe45LWC5rRyx0i0ynY1DxAzVzCrxxCOE/HZLzIJDaX6Jc4Bgdk+2
xp5a9+BPWk2MBGmyTnkm3EMsuJRNCDl/bekRcEkv4HPTMdCI7uhzwqQw7EAua44/MDiS9JTUU2Vr
rzbukTU9EOjVsqnBo5ji5DTMWwXBBMgmMXYpMgb43bmiaDmBTUYNKZnfF4ZWTlt5m7oolbsM2Sjz
BnPxErBbJewLOLA8+0FJU30WynxVw9AQo3vwo+/YRq+h/IYrBUoTbsyjy1xdD0eg8jeDXbWZmn1o
qf/yqj2KDqq5NwfhX6zCwfyIeFweLcsUa8E9e/UNfecEOaTJ7E26rBRMN0y1V7DfA6cVNew3KIxQ
wJ8QDKysTTVLoohs/kpqzmXhAICpFQ/JQebzZKjAwAsXfD15FuCjlg/XziKwacfcaVehSinLr4wb
Fh8JFSvZJvumNS1TsYdOJrkP8RNd6avEXKyLRq92OnAQoSiKuSkYVEydpEkE4rfdd26eXsU/8Ki/
WcMyRgEzCOwZW4c9OqZCYUFdxxOCRXxfRx/NgH4INt2N5M9D4UcgI2Nf8miKRUfbpb40C0tcw9Hw
eBxHH5wsRclB16MVc+9Svcpc79tnt6xi+Mc4BC7fkD0W2vurA5KE4wsWEGCbxfM5iwS5mLxgqHUH
yK2cK0tPld1ck0YNn8dYnZhl4EhY1oeUmWmN4fZXHnYUtpkl6YSEN06CfDP64oNg0YwfOr3BMPxZ
dJDks9v4i3xFamq6sgo/oLS9tRoi2U6O6nmfXN4pAPxF6Xbt/PwSDXa9aFa3uReM9K0PuxxQR+k/
Tem6Uak3r03qpSgrNVoHuLoT776I28RDqoJuFTBo++wtA+eHSeBsujQWbzayaJceZ0hMGMu0n2FN
6Pb2cTz525ypOV+lnU735/IVF7aaiw5OQjf7wGr9AB6L3rPbgUHoNipyBYtBZERAQH9mAVrI7EPr
EcMIBxG24At0FsCJd0d8DQvjO5r+3aaOBCFr+mEnYtbT2oLCmTJeSoZFdPN2+w8e5+pNmTQKNb5N
FE5rrbtwJFXeX0sh6biowwOOIUbHJEIqenO9mJD2w4VSo6NqJAPRvJAKMdE2eHrwMqt4tbduIXvP
AF5A6F9XT71b6lpfH7UCMoQvZtrKGONtWlBoSRf9iEjQamB2v+U/9sI9LEOiYH8oJ7yWpQEHrhOL
XieG1JPvkU5GP4V/ITsoFBt8V1zoEd1+7MM+OcBUYoOJv2k3lskjtFbt2CV5DHsCtGj6mjFT/eeV
UFKrlcopxvihwDGpwpzvBHxxaHVR5OWFOxa2sWDaphXrptqCHTfSpuGuQdrrG1f+RCye97RpVDRQ
3t4chy2EymvJdQjCa7WafT4eypywdGTCmeRjHcQvX5IOSSGaN0hnRHndBxXmmFoNPkKqvcVTybJJ
7xheFnX9Q4aN0Dcm1Wv7sKAftxmFq1zhRTUscnnRq3/ET2dpnpgwimNYcmUih7aQm51h6Bb/67BA
vlGUCnR1CM/DIV1a2lDgKN+gE1XduAaLo65Ee1rsnDhqjM5NZbTOCYoPbNWTaPgsoxu6X+bFIs1d
MGiX2ZeuINfa19UtoNSwYt68TP8P3Wc+4zWqoOITaV47waB2UWsPettBC8qhakgnfbUlO2/UuGJ3
1G4riylLvhb2GhaHe/0tLT04LxVTHiFVeeF1984FHlwgixlcVZpalZPhGHIvVxcbNUUeIDyVwe4t
fHZyurNZlVeuWcRqgv+QC3ZBL0LcA32fWW74C1NaXBSstjye4p+NEzz2SW7RnNvGcWIlbVRgjRMo
8Hh0q5b4VBHe78j2+cHAF/WCd36PQpo1eXi1HCuxI13Nf72zlzquGeIxSCBOdFtCA04+EOkPYrz5
UrvVtiuQpmQWXDpPrZcXXIm9XozKOItfeK6Qr/m42yt4uyoGKHWxRbwWGTRUP4YWY8DW/U90gfGq
vULt0p20ukNIucgkiXFLrB1zWfvOcRbvwCzRVHBaHdqrKEovhU2u78/fmlpc/rYsQEY0v4gH6GzY
0juVpX43L1lrM71lnuXgKNHPP08LQJ/FjTW5ZCClT2fbAofPMLwTmQndMrZuWnLAoVp5/gL2Ycg4
Tg3wuDAnTvmfIat1+xN0VDZwybltjrfPATQ7ebX0+7+WUbIx/Uoeaz7EuWi6p0AddiPpMLPCeq8L
4nGCBceskGldU7H6PCY7gqs4VzO+yVZteEKkJybv4XHag7iLDkSkGg1bgkeq0+3vMF0yvoho200t
76Y3HfmFJu48UOq6IVQG69Pqp/tyL4Z94P66Hm5tzg3N+j6SKZsIMJ0X1MUF5IQGfL2rOr/EokVd
X9kOyn836Qg+DiUN+7NZf83Qjd9uS+rvd65udnyvj1f/cuLYy4Kiz/szkK/XBMrba34xetU4+Ijl
dmNGMKgKDQSQacl22ldZneZlv64vF1Jx+JqvrfCdpzkbyOh/5ugGzlRl0ZDVkT3Q9GspWfdkmhtf
DpuoNncEn9I9xJ6RXJqnCQ5dLJ2HNDKlVZY2390r2n6DpSTWxqF0VrF4/sC6wnjkvMiU6o1JwrDH
wlFtcIf2nJmFYZbB6ZvDkvAlsZIv9upr8ctZ4zqmKyp2CLk3Yj7mida03wTIjZzFVvSgig45LSW/
yP2NxLQvQ0S4cUEuC112rOTm1YUHpqVPQSRVWD8+/ODgKqEwFkyCjfPDp57ZWtOPh7pb41CGMlMV
64/fd6Mdu+JPRmMpw5NbErwRhJk7zKhy9J9Mmy8CEKFFNBqSXunZdlrS/4myBEr0tUFGqi+uRsDr
lQ8dXyB+RI3ELuT7mY2vpde5uM3mKYAk4gzp9F1LgRfApGMLCWThxYRt+wMfC7iBgQhRPreq640/
wkmeDuLp5G6rS4FiYJIC+ijNQrc0ZJ97genZDvJ56tjRUiuEMrdIzsqJXsSkI9BZKVrdclRVCcqV
UAwdOc2mvem8Z5kD/u2+TnTDVj8o+Fuqp0j3Mc+zQeEHAt7cCvPt8voeZ+qsiTgFNO/OJh7a3Cwa
NoJjw/EWdCS3TOqGFNqQkK4y2rFCTzT3p9gAhMtr7phLFXMxLC88YbUE0vfgSjdE14CaIyKSfHvU
YZABMST85hynSu9rFMzKXMIwa4s4ELtTLRpcMng70VuegULENlP/nSD0fTRNVzT9yTc9xHi0rYkr
4ObGM7LISe5r7RocxhdJ9hUexdX8fqJZ9SqkFwBDLz8I3b+gUbHGIpzaaDT2qhiOvkn1MgipCuFg
7l8ZjjwPN4w81QXNHGIFIp0IvNmNVxUYnECC6+z/5Vn1rMoKQ1XcPfwXDveBAkAn/I6n0q3D3wGp
sZtk2ifS37I7b7iFmVVAhoeBYvC1UWTiONE0WvD1v42dshe25dhibCdxEm3rdaTK490ojLULMcJ7
vDgzrk1RqH535YgvbkGAE+Ob9vt4O8Nm9uMQB22CvTZ7FNRiJMefeBUXAKlnFwBMcd3Tv2zD8Td9
JLOBwjyjtce6renD51LkR8dg6tW2KG1m+YhTJFWIiOiXFx1Kbtq6c7TcLUsP5Z2R0/EHVLF9XmnT
2bjb2rew6yXuNQIJtNZcsLJBrUgQ5vh2Bl9rgFQNYjtjlH3/1qHSucATNo8z5vG4PIq3AdhU0kVW
3dDIMk0S11OYRpmMZSlCcze0RTgwzHxZcQH3Y010xlnPR4Wv4emWNEJhRAHPCJeU/HEeU0VWTedL
4MBHBQnyz0bKhNnLoWHXxHJ7exBFfmHdqEIfq6cuoBhqAaxWpjCMzLX2hGgknrdO2bYzDjRyyuOv
obQXw1VcWNP4pGIlpeDLrk/7CZiNX+zICL+rpPT/OXtNZyrfQn/zu3AFsn306ceNTX6Zo568jUk2
dPglD+csbuncf5uvotDBq0bMv4rsm5GYqxmFLeL59TT5QG3bzBfDQHgVSFwjMeMnZICZHCzXXHAO
J35/bN+apH5a3r85m83kZJMAj4Dr1rsWszrDAp7N6DxkbREG/JW+vkRSQJyUotNxy3bY2pOrxNOa
iLDsgJuyFzAs2C5yuq1um5ijCtOHbaCOYyhapAmoj96Np7G38HiHIcR+Fskh/KE5ibQrlFXbJhKQ
HAEMLGZYOzyP/yTGNTveTfJOE1aAFnxIiGGwyBUenxm1HXo7KzQ7kXpPss1Ffne/zTMIK+g0B4jU
QYtxo+2/MCmCNDSsozVrwFptTAySzOp5fEUdvD7zS7KQE98e/4ycR0wvk6EEFfP9/xt0g7fsYJzw
gBIcUF3/9LjSDw9x9VYMhinyqlqo7ZuqoI8C9ISGukO6g5WwEIJ+P/Z+HhVBK31d0Gwi+ZuIOo5+
FaopBIJ3yZe7MZot+oBDZviEfq3WiDdESpFTXEYkwPQiaGiWdfppFmtaTfhcaSUxfMyxL9zyhrPy
8HQLoHll+PSYWbsMfpER7UFe39pL3YBay050XvXzaaaXa+OzPw7GfGPpMJOJIOAb/c/5bditiJ2W
/qfNxhA5lX42BUrON65pAUAo124eCKKGt4ocd/G8n3STDHsA/OaEGptniFPagS9sNZC9Bes0/wQ7
W0VweiaiUHsy6Ge0g1ZfB9FnU4O73nr5pnk+YKgsqzIYG4FHAe7vNTNdVqcakZ3Q+gf+DgUE5bP4
7lT5vKZa45ZM/dv5QkV2kijuwETWvXqxreGhxhFGCLvXBFeNC4k2bW75diug22KES4OEC71eevy+
7z16u2seAmq86o7KzzsldZHmS6BFMsrDB7KDnUG5u+nW3xSP5zJgChSDemZYm8Z0WdkUNQJCVXDh
VlEw4XGzOqU/7U0YN1m2DqmCuZsRyqBMJeJtS7mczOxhVOfwDAuXpQZMoK43sCeTeA31Tqc8kDH/
lyrhLaClqTNUwbBJahf6Qdx4kZUL8+zT4ZDbIeanyVz/JVM4UrkRmpo4NDlsDvgZRcsTXC1848DG
OLLiO35n103GTiov0Pc5ktKE04G6xMr6rXb5u2ZUl+CcHE9iS8FoIoEJBDTDBL1//YNTwQ3SEdT+
LSaHqm7E7n1dcDJGjrRMPdPf/vOrkOF7ANALe1zNYVV4OTYzIjmRvUnVSuXFplfrEeTLPvjzMDMw
fkYXv/6ytSFBPXl2+z/tRbMO7HbxZrJlt4yn0Gf+iouG16auASOUkSsQDOp+3ids8YCjVBfJSwMB
5jwAoeyStDouWWYUFYKqI7g7nEJymI8KJ7GxvUrxb4NMyNSMdeVnhKOdUK5gY+BfKE7GifvdFwuj
Z6HymwVBkkM1wsjhHPK8WPM+4UAG4c+Tc1jHlMs8uBgnXrgmvDk44lQC8TFO/D88Oj3dITnoz/tw
YEVHu5NdDG/KaViwgH1eH4saLZc2yNBXjqtdyv46XvIFSyuAlMwWHoPVmEPYlS3L8JrVCYQkC9Ia
GVoeyCNtBarXwNtmHmSqGNYbhdb8UqfR8pDmQyUvMjrBAZZVhjtUJBdYq9/irjAI4jfleAC514A2
PSDFsYv9K2d8yFAUAWPGDIIlL1wVPA7pgkY7lWD0tDA9la1C+2fnsUppeQ+JHlv3HLWh0f9mXyyp
cKEBKpEOFIdc9g+FqRp3IYagjZqsOvtkxNhGGA/yLLKyJlsQQs+mOCT8To4jRyaxlwOui4lVAUZJ
0DIvKmqBkJpXKMvsAoAiMmBE8T14wwk/JgRsDtqFuzqmBTYNYA/v4uRau56PzO6Lus9sSwPeFErS
Vo420nQqmw3E+jhKxxMEw1Vg9XOErecmhxcecyzbDhwosbrWBXTUEIeeppIC7df9a/74npGFjmML
ZnBDm9zEWfCxf+YjjGkuFUk7J6Jxb1BpTYK26TYiKJporOnIALPJirDTGrjnIR5AavulD5BbEOl1
YJfRQvT2wUeBq10GTvtJwMVB8FNwatwhAFAcXuMlYX455tDC/b/WA3+KBQXKwklJPIoIs2WuXpTE
j0p5kkVLG8+Sem/RSrp77/GpbrHmh6Q5FdevRgMX3r/ZErlIpfWE5oNDUmiJvjOS/6FckCpvM0eM
KM52uWyF+kCOs2GVtPfznPXQkGFYdlqIQwRo0TXMWYljsAOX3rwSmE0aw+r4Efgpbo24a8qIlvil
ej7Osmueanz6KwXj+hD2hlKlnwh8YHHDIO3fcCl0dU8HJe5o94oB3hZ1RyNWW8pY4m9ZdikvRCf8
I4nT/Dbo7a6+ZlUqhA1p4mk7pCq7C9UjQGULmQJEilG5AftngSHH1WnkaIKDwpqy4SbuGwYaOitU
5RPuUU4lmAPMaBEogBaygYwdcvEOk+mDygOxQSkZOKTfg/GHdTUw4I1uE0pYBSO3UNniGa6tnvge
fDEdT258I9EjG7LGXUMXu4Kazajx+uXU06PrCFESQ2TYcWvau3yHaBiw8JiAYgvcZ9X5Ivv75emA
cTjgVastS89A8rX5bdjAtEuYUWQF4f7nSBT4EgV3TGM0pho/o7TUDq8TiIk56arM9fV5XSSR1lPd
DOvP/VgWzG3CWDrBApKZXn3A7FRPZIdu8GH9aQTzGMHm5mUFuH1yIEjFNjxYulMDZfroKQg7x1Ze
KpmoGV2lkgz9h96Treaa9jJ0yC42GLrGzdFYq1OhEnEkVMdFIZ8uYwSbk8KTqR4ZmxnafmRrlMVL
peSH8vS0jPz5t6Kn4efUwPTATBJniLyTkjFMEfKQsZQCSHALgUOMPwRMVG1zLx3B2EtYnpFXLj7a
ccQJ3fC0KcVcueFRCZP3eBnjBoOh2GzI897U9lp0ivm3Nm5u4SuPPDUEU7qU5tOCisnMqLrzBTYL
RwJPqD2HmdSA6JAIXAyVph7CL2G6gY0VNmoNMO16UlLxhuCJ9UYY9VnH4vvhNjO2Gc8sqpHWu9n3
z5vflu0tBux6aTFjpxoN3K6/9u4iOuX6cwHZjyl9/nR9HGpedJ1wg9uEpZ5XtyiLDf8fcQSxbG5P
LoybZbN0UIS+rjSMWClj89loCRtlpTQbn57CWqHDaXVq4KV1+6R2Et/4KXFnqB3w32Y5FF4w7SfJ
0Q7x/KJZYsdEfkXHp2SNdt48vYF/g9qNVnCg1r30tVoQkQVBBkh/vnuPLevL+FnYcpgAhtw7+vhj
cMMog/5PWZnEvSEBQ0Y0PKupY/u9EOnF2Ngmu1ldpbdyKinogyfBShRVAGpiUK+VlqlZIWC9gSOb
O7gwPpJgdW1DsUhwf3AaYEU6Jl6WnpOQlC5FhPzHoLHkmednFKnwkhCYRwa2qa76KRMp/ymAwUyJ
WLu1xPXfKy2ZBdnnVUtgQPFU0eOnpE40nzRhnZc8wX0Cz3dzz2jR8oWEndDcTN16S8HgTDvzflI7
/URYN3tGeDnC37oRLj5bPe0jYxyoBtJV85UIe0Pq8lDxkmjUC5rKJf783vBNRBTBjtnlCCyDjrym
xGNpTTUbXXrg9NllJrR9+D2XRAW2U5woAmHIFdwHep/JbA9LR7QCTfvp4yHHGvcAvIf1N9oBf3QU
7CD9BBtEFyhRMWVqPVyGOz7M4vscQzbbHlNsx7qDFDVqxv3r1mEpd5GDsgdLZHRGKg9VOnnfhHMa
qmSZDJidheA7fq099mNd683EIrjqVlE0ewMcqXM+0eowrrbHGxOg1oPf7orRYY38A6irMXxfXueO
x2IRPkUGmNWuI9xXClZfR9VJs9XwmjOWDJsRZehmoQ/wHFQ4rbogW+D8VQ1pKYd1FxeJcCSfLzsl
Fz/1Qq6o+8iWD8C71Fjui5oxIV57cL6zajHFLtlIR2w5n7J+BGLoMWRmulKMclL8x7VKJAZD8yAt
Xt+ypK8xn/zq7IcVNP52CBbFNHt82bwiK43LfAMa+rb08QWF/sxeUGXuDB1xwOOyequfXo+4smoR
KF+kQGOMSpR2p+hPQJ/GTIWPbtY45p6lihhaLaNmOuaxRPi1aGthE3UqR4sNM0Y/oxrV9RukhMc8
kiqUsjdI87wwFqDSdz4C9FaPwGKfuv9t0n6thOAzvqozHaaiLuAjwxuv3WRQsDLQL8yhRhNgpmSn
1UwIt0HLNxgZZy6Ls1TEgb4/y3wIIYGxFUaS691w0EukhDLztxECjSXidygWRpuz8cprbiQ8KxED
OL453vdvcJHrRjSlYsKES0F6K7Y1aav/7OGb1YTFSdOonXZcdwge6V3h8efmfAtEXc8YAOVL/TsF
ls86IpPVIljSLYE/R9Xf9x24sHf6q7COYzlw7Krhl4vKaUDl+cIyqNqMJTIix8emddl4zUwiF1Rx
NRlcCNdr0ZAPJwckLEMGZ1pj+t8Pbnbh8qbOi0ShRoJ1h8E1md2JyydqA4oo9qzSnd+Q8Q6rK+jY
3QDNvtxwg2gY0aAUReBurV55ZwnSBzEekd1gEukrm4RZz5GGzqSQzMyq/IiZCoK6zg7NTW/lY+G7
CyJtUc4OHi8yD9vONb3wSJfUdmnU2ZvT9Z4lHxiarN2+AgQUbraXbzGmQrhMFo53AXyDspXqTWCO
ZhlJjBqnuV5m9XLDWLr3e/670/t8eXrRuYhhZbKnUmRLdiqNWz9w0dFEQIqdKr9n3UI8yRotAd7U
WDr7HYj90JEXV+xhPzUO9HzaVPC9K0Pttz/FnMU4H94PpRBAMfWsLvd1P/1m4ncMOxEAuBUuz7yw
Iduu74K7AH23A9qun8TskYQZ9lRczhPAeTwmlXeH70GxOwDMdQ3ACLP49ropFxnMGHdqs3SFMIWu
0AxKkQDNbfVodtFXVS1PZP0X+ZOIPWd1xasieitsJ2948geVFTOYJ+lm199TECRroXZEHmVlFMPA
q+3qAIQdLuyLMg/OLVDB7kW3KfX2Zw6fjX61z5jSYZRG3xgHiL+Qlkx+sPP6fz2yqIlMHGn/lIFl
NndoGeeGNfJnpyK+hCXxTo+Opg1bnrgJPmC9ZCelMZTMiqtpyhSSDOyRbKYWahbJGnh+FWE/aHV2
ic9hUA7uxTT9Z29beStNVVF9CUbJ8d0IrQH8x5kGMnXlvSYrbCpHvhM1KKzcVRkCKUgJYsqZvBKW
HchhyjMgcpWtWYowrB7AcvoLhLxOIb02X6BImHWF7kGp9VzttgAAvJ31AUUN7x32+yc0RiVKZcsh
DKqsPRDmBesB8vZAhl35mMqCx26/9EY4ywdREr6xaziblYZUT6/KVHpHYAacW6o/ktrONbrV8GRD
4YjWQj2iJGi8TT/jUsloOw89NguHHuseUJBkJvZ7KepWzMEHAVFVcdkQB4OiR1bW/BPYo9oD9mI1
VZAy+i/tUeqqcfYonHxJ/DXyBLC0lTuNfG7oSVMbY//x64wACOLaq1noEoR4RdIylQ++II/AxeQg
6Vs3rKxTIVOmLazGnr6xcqRrJ/RMoPKQNIeHd1aFc6jUasZZEyOTKWQ/7X5xBCt/ZpXKJowz9e/y
Fh8TVZBYM6Zq+hmhiK8pq+opi1PDE3yHJTr/v+GOYa7hKVPZFo9s48fWmEaQQCFGhk1DNAgT6tw9
gR6awwLzOxIN32BvZ6Vt0gJy0iCMhmoDQeU4p+e53iafaH9GRUhYQEu03RnsUvXtMLu0pdRz7gER
Vy6tOgkMdd5DXN/z//SaSTOuoCE1aPTCt2dyypTxLS/zBSmPPqlJ/zg1MRy+P7TOEdh1aRS4ZWyr
nDzo9+8BpDKCkBdWbhGJG66DSHW+9bJrlzqdTJ+0VGD/cBsJiXDrNvkgSO+7uJcAQw+1VOMGBIal
SIsv/KXFMQ5ZAnylDL8wguC31EvpAMKj+FbYu00+XpUoQ2lbq7lA4utvFPdn/DQhBWFVoZxqHTJZ
qGkZ2+UycZzcKCdW7rB/guerFcboJ1A7I36MB+CTtSEL+PQJJdttzjeODjErxP5kk8VsD7xUnFZG
aj57HoOaa5i3ZyLgFSGri8t5KwaZ+hQHX31ReAC1A6NoNU29nDvvu0NsdoAE9Y3ZTtj2ws1j5FH+
ikMV49jVWD9FBEUtB/vcE3g+ZdWOzNYslVPyDYAqCOAin8oXUkOUKHP6r1mfJG5rdQEDGMTdgjd7
yOfWUdQUYfVvtr6k/8rY9O3fubBUsSMHKFttUA31KKnPJzHioi1qOTOzg1V+ANhpoaiCsJquFIwX
0o/kGeevoy832R/MCfK5oRq4CM/KzEBp2LN3arUyNTIhEO9epLQOWAGXF7XPqjMpPbyUAm4U9S5X
DcKJti2sK1pPLo8y+OvtHFGwNl6SVFup2zclbdDsp384kN6cVa/q+2tdp3Z4cMRtfzSDMNvL9x3Z
J8fCPitNDEweTQIOAtXPwtMzoXnL+4pn+YIAKXO6jrm96GmxQspGzykG7S6IwZqMU5v8wQ1N8IIZ
lRImKZGPI81+00uhYYStSuxB+4hZSxpK8O3zPtjPaaWAGqxaaJdn+A3w7GP8fUiFKjSKGoWl9UOL
4ThMhFLYOPP2yuVBdH1NyS46JhJfCpWAUM/0SJcrikZjH6kt7v1lll1Up+TgNfXO7P/ZZaSzwsyH
fvaKuKRedNVjKDm905QbHeLbktAWen1mmXwlj8+6VLwGtIqb8OXyoqBSxCu71covWpb4LqZPRWiC
qsFuZF2109ogqtj50sKAlO4VFk3ctg0qeHaDVezAw/LPWZ6PAqxxrXc0iQIXeJeb5FOjPgwESO3m
iZb23PYYgKYghYc3IWd1R0vbqIzawQUaBZb64uzQKeel4n6+YCbk52V4b31FMmUP7b90N1Ej4nRv
dh71XuIKawQkYLAplOhsX7Srw6sBQdZQlutiGx6tHq0i75sysjXN/Cb4J/K1zGwFNAei+uHLae8Y
Ghc5bFFQKkO91EEAKaFWbNjpxDrvg8o1UJm+aHYo0jrfphK3sygatwJnIvE0mk5SBPlyX4EAK+V3
6egVsYZFuLOTGoK4YK0QtwyH7IEGVklwlFFvo4n6myPWkbJtStYiOvAkukDlTHsnf6rKzT+NzxqA
UW+2CC6aG+ogYb77pwuu47yz1MRAmpcgOnd9M2LnaOY5b28wHfFpUj0ZpjFjtCJUOMe79uS0oaVJ
buj2O8d+VGnOoOmc1FOwt9GnWJQfz+FKpkDLj+j4Gw8ZlqHashTTZV6iNEUJT8xdtctd6oNk0dD7
iTWO+YsktDrYKlEo9fcAtrXh9RcnkyfU1fP7LNHrdObmxNC7i39Np2fU6GooHpGFrBaZvbTrzv8J
CbN8W6NgD5qRIoGJu/EKOlGP7jkxo/tglkBeUmKpUdmdXH1+EiqJW4ReA1P1TLT6QH1VL7ELLQLH
7JthjHRntCdLcEv8EdFFL0xBwGUPx/waT4t6mpzWltCjEILzjOjlHJAFbB2dzeUmx1hpDVd9JK9o
h452uBfWa7LZ+qG+RO0H94wSRhmoN5lcBIhOKrdPfDHYgpdo20TNr4sTQNcYuPUlxJLckatbxY9n
KxoJZ6WrRxgcqeSkZEgY8BIkbLsLwx+T0w3bvmtgjcIOYIzf2KQ4/y7+zTayoiAvBeSUgCE8+TPW
t/gJGOQQbOJ1Rd7xSjdnvvVbL8q2wtk5peI/hRwV3cTuUSy/d1oLyk5BOgSa1BZ/+sfaBVEhSkQF
Jpj/ayD7965Urv9BETt28F0F6R6RNIJajhmsEZUyi+Q0gx0RQ2K0lHjsi1GfTEgkfddFkcS7c7Po
BD3LrMs84Iw+4SiUyYB8pUWqJVxNhoOWOCqOW0d3zkwbXUQQoBcLCNARAqmx2i1/ackOB8wcUvf9
F8aSxLKld3JZKYfaTKXtIQe7xVq/P0EAPS+hhy0ttfRDSuLFY6r4KpiHObUVIyhrTNM7a4eJS3OL
g1GYXMcY/hTk11WZ5na+iaYnLZqrg2QVRvGL1GuEDO2MLXxnbdJ4+zpHscFQ0KZwBLUACvK0l/RJ
GvtWhqpL3xfhbNc293niS7svmAZS1tYIwIzQNYbk2q/PsIdf40qucQPwmLXcqmTxXa9gBY8min5u
7LDxTawJoE4jdkJM00t6tdNw+dujMuWNsy32oVt4NkMnvpPLtBtUHQ51kIxnE+mHvC5UqAo83z3l
TbfDvOqinx3NEaZZglIGTOzRyFsLzplnd8in2dZU1IWe2Jxyv/bs9UbCfLcacnUIhYtrv+Dsu8Nk
aDonK7ivDqRKgHBEO9ThO3P44GOdgeH0To8S9CeJwC/XvCgBIxVXgYXy5dSt8pqDosnTHIwq9E1N
PQgVYdEq9hpeQGSRrxAMs71CE1+N50Q74Osp9TE5+z/ZPKPTbL0upkaND0p+Q6jk/+aAzEcvmK33
FeOULPllCdV1r5NKMYzeBqatB/me7fysVnm2GftWK4SzIiuwpaflGAw1b8J5zRhTgiwXaHOmUL5w
NQBTCiYOm7mPBDW2WE17p9t20zrN+3KyOU8WnXQr9t7oL3XNxjQFoLxiRcvIp5iknZ2H51uWaHXk
VHwEVzFHuhwavtLul4oFKm+QICMb2FF1fv1+9MOoH2HnDttQUxjqhb4iILhGaVEZ1Dj7CczF8l8t
Mjcd9I71QpYFGZ0B3EjPuI4O5EdjCDESDw4sGazadqzxUjgla8cslNfTRwF+ctytgx1kl/y5IBRD
VuGMpg==
`protect end_protected
