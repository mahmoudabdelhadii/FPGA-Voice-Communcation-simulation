��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����N~@#�k�0!����+��=L���0�ԴZ�2�Mc���ZO�����=�����վ�	"cqw��a��TS[��{=:�����K��-�մ�(��k��N�-� 偙O��QZ��~rL'�x[�i,mׇp���O�I43��4d�,�H�����SN��d���3���r��m���̨T�I;uj2Y� Er�*p�Q$Gm���p�V�`�2^���,hz�<p��l�Bxt�5��s��\yq���#�@W���f:m��T�	,*�񞭋����_��㧋l�	�\�:��uGd��PǷ��N�I��_����Tuv� ���us�(H�~�{2H�:Zor�Q	#%�3ˠ!��iS��95�,?�.���/�F�i{#���Tp5����Ҥ0{%���2vpn���X�����@l����3dc�ק�3	�Ed&3�ZN O���z��s�yxӡt��v*}ԫy nj#��lc��m戭k[��5)�A#�����8�!�]�Z�s�M���t��w�!��'ÒE�rv��Ϝ�c@<U��\tq+��&|�&X1)C�����r�A~��B�&�����s�:n{p��͠R�X⺂L^��R����c���f��J^?��ܣR�O 1�rV���:��T�4���AD����˩�F�w��)Dm�O�b,�a���1$��c��7t[i2>�ޔ0,S���󧇳Ϟ�ᒨ�-��}�!6��Jyv�醊�^_�(�H�(y^����o#����X��3-�k\8�M�T�"`R�DF6ȕ� �,5�;Ҭ C�k���1\������k�t־9�}���� ���QHF��"��t�9 ?��{E_�7��!����]k�j*�Q��~�=�0z����o<���_TC?�];iW��M������O���R�$�lIlqֿT����N�B���ڊΑ��R���s5��yEK@aTaz�]���@	Ɔ������)ɏ�������7~v����}DE����S
�|�v@L��_.؉7Kn���Y��?j�,/4��X_�~��ڵ�W��S@d�|s�(c�8@k�@/R��vk�,l����*���ٓz_��
�
 �+����]��^�,�+H�	��zF����"�~i�Qyy�K�LR�-$'<1d�X�]@��N,yی' c���	�rݒ�$���#Im?
��I(���Fqc��g���׌�]>rgQ�ĳ3�` c�	\�آޣf�`=�C����Ӓ�Le�͌����aD�8>^z�+�����Y$����!���Y�W�s3J
�ث'��� �wJ�%�,���S
����)9
��Im�"�PR����MnY���"�{�#����pJCѳr���^wT�������f���Uܲ{���E)��f��wk��!�*nn���k�*^�	j��;�S���lMV��j`JՋ�A���G_�΃������A	f�F��h�Dqn9'��7<H.��Ըo7]�L��j��{��Z��|u�#�ˈ�[+�� VolJP����]���`\|*l�2I����<�e��K\�AG�M�7O�U{0�]�@o�}�sO9�5^9�mԧ�e+8;LY}�i��N��0����Ϛ�7#�.����v;F9bn�?hЙ��O�.vBgJ�1o�(5��7�B��V����ծ���h���gǃ�Q��/��N׼P�$��W("�41�� ����3���o.9��wST����J��*�܂ꈹJ�	��i����^������.a�\�Ǜ*N텪]d��7�c�j��k�����\J]�ؙ�=o�J{�����(�os[Je����ɑQ�E4W��	�	kr���Y��1�F���_M5�no�g���abq�����ߕ�(�6��Dp��a��a����n��*ϛ�=p������s�#�sb*��C↔EjNJ���K{����e��c�_�s��
���i�y/�޹)J�dEV��?rjA����FN���巩W��D���~��2fT����Ug��{�-�ZZ��rb=���aD6��A
������|�{�c�R&'t�T4:���}o-���S���f�O�.��G�8kBc��V)_6��4Y%�O<�
<�(*�'W%-�O��EI�?�5���5�س��%�~���?Pk�� gm��\�5x�����ڐb5"^��U��2\��a7�n��������b�3s��s.r�2�M ��r�r
�]gx�]���>�D�&�\`x����Ra:�L��V���_q+��g�IS;��{5G�W�̥���\ė�Xᥗ�U!����<O���3&zjit�K�Q�
jVm�Ra\6\ڛ�PE�����I�iգ�+.�&/���P1-�QO�󠌈p�08��*'V/FO0�����+�X�kӖb4�����]\���_o���mI��\��H�&"'P���z���jD�v،us���e8�B��"�^Ǖ�Dҋ1��M���]�����yl\]�K�{`[,u'����Ƒ�
y+��Ft�����A�'��D�*z�?�)��p��ixZ\WI3��q����G�3��''��W�[�k��������5��%)*��x�۪�f�绍S�V��r�(�\k��K�E�����ó�z�5�!��X��I�喩�sR��Bn��.��h͙���X�,w8dU�و6��LH�P���"���ѽ����5QdM���]�Ӓq(��A�Zޢ�ӀO���Jۇ�W��q#������k2/��}�v	���!uӡ4��AM[���7S�l<�.���O8̌0<b�r�h#z������4��htꁞ��7��Ar%�>�K��̀�v�S�=kK5���.���9��7F�c���L��Q�N�E��z�o�鰢�.��nD����D�`�9�߲*T�t������;poy��a����Dt��5�Zc���_U9� Q����PK��5ΖD2h�)�[FXƙ뉪��	��b��w�D�[�a�ۛߓ��Z���O���,אդc���EC4�ɕͦ�%��M�K2�E�^�g;�)���y�N�������:)�T$�A��h~��F�o@F�h��E����1"�r�T&+3�"���Ɵ} 6XE����:꣖4O��5�إV��M;=�8H��:?	A������Lݝ��,k\�j��OȬ7:~'s�5k[�gk���B�4o�Ǉn����1Ľ~�v�9b�}��5�зIYgk�h���bfw��[Vͼ(�I\�,p��@d�}��,���Dj�	�y>I|�䋔(�8����Uo���?w�9�4�;��ч[f7�><?�q�Q�)p�����e�C���b;Tpn��� p��3u �d֢��e����}�P�m@��b?�Wu͒t�ۂW��ޗ��\�C�0[�J�{�q��J\N�L2�M�O菾s	]��� �}4�#b=,��Y��̊@9����jF�j��iD�T��ͶCK��mO�|D��
0��0��ög�t�c�.�m�1b��w��wR!¸��@�I���0鳗<+�����5>����j�P��/q9�,C�Ҥ:�`����HtU��X�.�ԝQ)�Ɓ��6d^cধ�{U��L;��XQ�1�/��܋(�i��!��o*lz��Lw8*�U\�)[S��d��)������|�pC���4�
+��m:sz#��{��SMoj���Ԏ4��@<��#a�zO&��^���x�:h���SP;ɘ,_xU�x���d���|W�+���T]��gs���j��� }�\�}S2���LPJ"���r�j^Q��i];5|Ҩȗx%ټ�BeMv���@���ͭ� Rm2���T�f#�y-ۗ�Wa���5�4t���V����Y�}��X��f�-+������n�<M{O864%��PV�A�� +^�,!���a��a��&�V� �D9�%n�?*$°\f\�3c����'𡒫�B{��
�<�>�H`�3Ǻ.�O�sR��ʣ�Q�[����A?�ً,�(_3_&������.p�����P\w�:yMN.�ФA+�a��8� iY�	q݂��V	�g��<���qP��70���+`g%A��n�<��WӢ&�Yh�e�[X?�*���	��Qɦ5���<�y	J�1߃ a�T�]�=iƀd����6%L*O�&̇���eпg��O�^�k��+vς]�Y��D�>��L�CUU&��&G������O��~��Ú"kO���� ��f�%��M����1L�B��h��� �0���Հ����gZ�ͯ��P_��F׉�'�0��yű�4f�`gB`�(���tڐ�5DU$ڿ�G�t�7.+u�׃uW�Z`�ad��-����Y��ä���d#�6�tpD��Hj+�v$�����B�T�ϔNK]*�2�����ZDgx{8y,� 5�ݖ�.���"lܯ[�AY�P#Ƅ�s�6��r?�Q��r]��3��c���@�D�vs?���e����������j�l�<:�-br �7�-���l7�Je��c�(b�6�$(r*Z�8����d*�ݿ-��A�Z
�^�|��U�jZ(�S��:P�� ^'�C�`u!��~��bu����;%�յ\F��=�o�$s-x�����גqZ���� <��ATptE����-�8�.�5R/��YE�QpWw\Pf9�����@���廕 ]���P�],D����POY���u2��&��60rG�!�3�0y�Y>#�⁵���%T
$Lt����{2��q�~-��~I��"%xMr[�	��zxk&�pW�fm|U����i.�������X�'����~��Y9z�r�������dL���X���4;��� 3��j��<��W{De3)}OV^.?n����I�&�le��	�f�����y�Y�<a��������o�ٝ"K90de����V�FX�RQ�a������]"䘛�G�Cr����)�C��NB ��"����YJ^��Tx���=%.4�{��G���:K2��ϯ��b�h+�z�.��>v|�cШo�gs
"�ߖ��|��#�q+v��n�d�2zGf)滺����zL�O[�_Y�f7��C	���z|f��Ӑ�oW�����I݆�ʿX_a�ta�J/m��#�)���K��G�{j����6Wi�vZF/�9!��:�zߎ��Z�)P4�ܦ�(H�cA�qk�x@�*����p����b+;B�"bZ�eA	��j���>���Dv3�_�P����������}�+{q2U��۰U֥W� ~t�<,�7������M��9=bTJ؁'@�ݭd9�=P�E�rk�|���T�8�l�������@�����H<�)�?|���>���+�����3�-�}ނҲ�T����:���2�0��l�s���'\�F/4@Q�nל)N�%Nk�M��d����n�\�:��B��t���W�6�V�8tl�ˎ6���G�n�Z�����:��^IB�P5�H�;�Mޑ�]����'a)� bn�|)�@�У@9��GE=ƫ }DO��>(Wh�y��hA���Ű�U�^�\�L���
Twh��d󷛱O�jMv*㼟��(�ɨ��\̟q; ㏕S� 1,��7���Rl���Dq�B;&7�Gfh�L�g���0n�TS�xD��N�O�Alx��'z�4ľ��BQH�g�����䎞��0���!�z�/�E�WQ���@l�f�dȳ���ŧ�yO�Z��s��8��m"s
wGZQB ����0b�\FBA�A��<����	��UE��I�f�Ñ��v�)�X�����=��j�I�,�B�I,�N\����Y��$���=r{AFT��˨�N�[�w:��)D���m��'-@�&W ��2؜�ٚ�oG��������AE��ۍh��8λx�ך=���\��Z(�t��DNêi��h
�N���L�I}"_4�~S�i�Dk��RM���]\�Y�Q��a-G�Fg�tWi`r�rp�l���Ř}.��x�c!�U�q��a�SZ���󻢇�̟<�r]���I(FB��U�q�i�j[�FI�M��0=�⊡*�*�5_�tR��nd�{=I�3���{ ^L�^����h�R��pð?-�&�3b�����*u��򰚰�n��O���^q�gjt;a����x����Sn"'�,����QH�g`G�\��Jbh��v����u� �od6k������]1m���` �k0\�ͻ�������L@�&=v0�@��&_p�������N�/��� !I��c�W
B)�����ȴ��CI��pX��|�
(���Y�� ���ޒ��*�1ms��o�,���-�y�#���o��a/���@7�r�	E��S��A#9�<��
֟��#o�	(����-5	܆2$>�
H�5V)�5�����c������V��Ԩd�64%|��(�2��!QA{m�����8�D+�S���8���B��|�KScߗ��=��Y��{���>�|�N���F���K����7�\�[UƏ:V���F[%�2;�[��n���驽RqmUX�,�M�K�:j���qP���^�Z�r:��{�%�y��=�h�o{I&�^6U�G�3/.)g&�4ƚc�%��w�BE8��|�Ͳg4�aץ�����*��1T6�IԯL��Uj���E�,6XAԷ����I"�g�����!(�8h|���_��,_X�NC"ˏ�%�)u4�kh/����fb'��ب~��U\aj�
�_IC���bȼ�����`�]J2�ɜf�UU[X��M�[�4�u�!I��i~8}���&'�-1t0hèc6/<כf�7_7˛F���p���LdaZ�$&���/���<�A�#���ͦ�*��� ����ƣf.��^Z�j�o$����Q&m]H����ζ���v>�wiϋj�tmG��9p2Iʆ?�ex���'��F/���V�
��=��S�-^M*s �0"{
������g��~{�8���$�1�7).��^��(@�'��ZH��]c��U@�� ,P-�	���2��m�>��.�'���+k��ɕ�<v���E��U���r]��
f�v����#��Rr{�R"�2@�G/�u#8�%�:�#���A&zF	�LL�a;����(����<�����K-�l�x>E�pKD�O0���ET=�ۈI�a��Ư@�qkT(�>�te���Qeg��e�]\�0��BH��15ki7z!���a��$�����/��òFZ!����Y�d`1�Iu�o��\hzL<n;".H�2hA��݂�YU_l��?�(�����˴�H���R"H���[��%�mQa���W�/�yk�06�����b��ܦ`�׍�<G=éb��>��Xے�|�
H.ujP�Z���YJ���w3���[��Yb]}������K���e	E�h�v·��X�SA��Y$��:��� hߩ�N�!S{��K�s.�!$(\#YR��m��~�'�&��"^X�c@&�\r��ps��VN����v�y�v�Vd���X�(��8-�W�`���L�5J�5v�OWH>���a�+2��������ʟF�2�:�?M�x:�r�o�?z�z�\y��#�s�^�w\�ܨ�?��Q�r �0�$��P,��95gT�{�G�n�@�3b�{��q������'sJ���CxIjLL��Lh���گw/�.bt�:��3dp|q@�H#����n�b]�����;Q���c!�����?�|@*8�7�}|@D��ʳyj$�N��f�R�z��p{x��^���&7%���.�(�����<D�r-���vw���j�R���/���is=���$�9U����"���\�fOdi�6]�̝�ܞm����9�m7�$){�W�s+!��F�
���n�{諦j��7L�'wX�*�-3�҈x�m:��ʑW�[�u�E�R���|y�CK�B����&zR��fl�8�����{��X�|���H�{bT*�%ů��0�.+��[��#�E"x� n �����K.^��M�{�4����g�����?��7C2)��I^�~Sh�QUi�}��L�M��d��/E<�=ޱ�!�^%�{��� E7�Z6n�'��ɕ�ICl+TU�6j9E�R�I�~����l!^)��N^����0K�ͳVa�M@C�|
0��NR<z�*/�Mc6�d���_�i�s�O��.WI�P��0j��'4^��U�T�����Oahs,�F��9��)E�gqqqK���I �����E)^rt��2L��a�0`
��Ŕ�t�Ȅ�*���Q/_��Zf����}�پ.G6}�9I
���[��a0F��X�7�h��;�l+�g	�T�t����!�a�"|��/t�1a�(	D�qT꠱7�}�I�R�a��?��*�RC��E�'3N�`%���ԞDib�ݢ(�ӏI�=%�6��:��{��Y�%�Z�����}�Gu}\���Ȗ��\�Q#K�ܪ�Wc�I�ʼKh�����n�L�8H�gTC�悈�%��Uu�*���5�����Z�4U��.Qq�<(~�;)&�^�gZ-��v�xa��b����č��~��^��1�\!y-���Yu�{u�-A�$I�]�t�$ wmã5<|�l9!p��Ԕ|�~�X=�mx]�4����H�O�����D�I�����Y\/Jh}�+t�w��~4!�wf*��U-Q_��+6�ܤ�Q�즌��(�����W�6�~�<�K#�lL��v
�G��7�ml��1-k"��L?�G�irF\����g���<�x����]ķ-�*S@|�J��~�؈N�[�+��+ӌ��N£Żl�'����x��L�O�5=����vN�ⳮ�U>�>�,���4�ߕU�1�d���Q�B�f7Xנ9�S�cv�@.���V=( ����*�G*�6��z�ߑ�Όn�O�dG x�3b@��8�VZdkuf�s�48q���C���C�'��P�q@,c�m@�O'��;SD�f�� ��Y��I:���a=� Z)d��7Y+>�Ӱ�~0ǉ��+��@���b��R���0ܡ�Jc('p��^�ؔik^�Gª�K#����':��u�C�����ϒ����C����й(!�{��@����j�(M�W����t��a4Ң`gϕJބ{yg���
bq�&y<q�2f��-��֨Y�{�u<]ٺ�@<_����P�ǆ݅ &	�M�pǍ��\�K�=3�sO�4�����hATJj�,�z�m�U���\qB��Q8��Ml��y�;����s���gw����Ӷ˨>��p`_)�4��m��yg>��N�f\���58�L��2yZiulv�I���<t�R>�A��L�Y/��⛚�������D���?���`8<ceHUo�'2o�0�	x���{U�F[�p���X3���9L��K����?����6k��ѻ*�D�����@��k9�.�2EP=������"2�bi~yd3�u�"-�h�~�s׾�8��Q_�Jc
P�RM��Jb�t �u�|���E2`�|�;��h�R�����H1ht�xp��O�H��}��B��T�#��Tի�圹-�����H��Y����C�#�l�8K�a(�¤����U�wX�8���Ot�,;�<�
�a���185�3���\��hP�a���>R�Y���f�Wb����+4cH�