-- (C) 2001-2016 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
J+XG8RKZvBOkLZtLq6PC4A2n4ubt1N8eAWgzjiZ05oVt5rujY1fGFoCw8UN/sDZFSOKL5yc7NnMr
MJL+WeDsixiFOjLkn/QdZDih75TbJdNKE+Eu+ct7BLkF2En92Css0Bdc1aKZumQ4+mNmjnaxzUU3
EPBV+7+VlaT5DMEGg10SGXN7+7xl4DyyR8DuLJENnrpYodyvBNWo2OlVN/hB+iESfcwrgXW8sz14
k7aMYy+EekSsVT2bJ9+w7f2a6NiNOOuP85LH+jRVu0Yb8q4QFRbkwr9+Oc1TKQhVtvnFtEs/DCZQ
8JKxjU7w+9dGoLTYBk3840c2aU7YSABX6wtTIg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 14848)
`protect data_block
7XexQpm2+1ohl988Io9cw53aJAXPCxtaEdovbzNLfO+yyStv4uU1mu10fjU2pokHI4hgZfBqxPNv
aInNP9xwhhFEJrsVPsaMotCXrXQQJCPs4OI+Mh2o0f4ONI22xmPJNBYjn7E6l059zCCNcVifXP64
2d+FaH1Uk5dfzPbhXoEA2ryw1W3chkuQLljsuJUK2tOJwymOHRG7E8dV8dktRFopQHXhsZgXKuM7
Yc6AzDQelk35wVWLAWVi3wl4WVhxY6/IR+nGvnGDqDgfpXRg0889XAjO7Xgzmpwga4MUnsMlMYwH
1MGLae/JKxjquynlpTGOcrmIv8hJNY9Ok4FkputNdRtR9ovFchuooNCPDBXR0l+1T0u11pLceqmB
dVFMjKPKv2LlCOeESeGvW2Gy7RiHpQf38LgTK0lQz5yRUMMGWgniWr7qMQsWq9zz6vvdRn9c/Zjy
5A7am3cdqNd4vgzHb7W+1UmQUGSvYQxxJXtIuGHjkU6nItXPgFV4rm1fGlQdHwdfGNFWBZWkDLMI
t25/Q2v8XNGOYJVlXo9D9YKbFI8C55MqKm7sD6P8pRGtWJKevyzYaz7ZU3gcOKPyOyTGncZMDoG4
cLUija6HMmFcGhHeeGygOrT92GicL6pPjgfeaTcmRmmH9Pt0WMHEbKf9ybY7P5cMqDNCYFn+zVnu
ysCRXICK33ACMLgTvPywGPTABA+OOwPQtpffaW5cXd1YixzKNymmKKDuThDMlA4IF7mc2PrAk/PL
BvtqGRHcy5qhQ7laeVCSOBWzcakobJKiGhcYSoRzpBnJlP4ibbwIx+2YrBRlu6kReEeTi3rXKKax
RCvKLsporSD/2EtKd1aADUQbS91Kn8FvZS4JljKhGRmHS365yKoSz91CCIguHLTOi7xa6Npst2mH
lQFcWng5FFGpEqXB35NdWD6FTt7xnT+pz5GNy370YdZGJw/MPNBnJNOQEI750UwUuC0cyP7D53YR
YgqPZ2+px4c/xKr5c/aPe767hb36k4HnoVwot81YkEfZMwFNbg7NP1VI2aIvFtJVmJuqsCDcY3+M
JCMhZzHlXuS5M6MWn0ZUeKAIUgnSrBheHOCTsbd5K6osvX9W6heITyWrTMm5T6sNgMuQn8wCj0Or
OvaQZAViF2RTsQbjGPfYIz7osgDBuQVaCbzy33FbDy9OpRiP13JX533M3kHvsPKjgNPauMPje17f
2hEXOigpone1zSLP5Sa++s2dEl4b4YM+NnytUpbI8FC9OM/Vt2PDSgPlVLmrdkFMSRGNXXxsC3oe
y6DRy9rX3W8r4DQ4xE56yArZP3I4ZYlq4Mw6/5ytkUnezBGIm+qCDpi2RLGOu8jIC9KhdIon1xWq
LqlGMAlCLNLCn/pdyitG6QWmhQnhepSheaD8ZrxnuYdLac7OS49zVhlXI7dzfEws03XTYX18sYWn
vvBwYBNeULNijqpqmaGQXkauzqE3fnN7v8us2KHsTcTQ0e613yxOI5qrHY91IVNbdUmRZbyyhtLH
P/eyEAGpedQuZCw/RaIujHC2eIDLoWaP/lPqlESudgyfvhoSXG0uo7kkLQdqYKIHYAPA4XVJtpxX
zGKEW4JlcE/xnCHuD6QqFEQyFUj+ZwrSH8oNfTz9/D8xwr9wM70Ntp6oit2/xaw5Cr7kEGxm0KBW
iSs7guwR7hDjUSbZUKmMlDeI6wwJgVeQNkIK55dzIze3Cdb0BtkdDbsypP4GeULvoMj0+Z1OLKPk
IWivrCnl2s6NWSwqokecjJBghDJy+sxd0qyC9Ji0aVsrnp+toQl4xvq73WFyppxDP0q4w1v/ainZ
+7UyoPdl4mF7JYd/DqEhZP84mtbIXU6+sPSiQSEWA+YP8s2soqSu7cqpE8s3i7wvIrX0Mizzpp/v
OXFkrRPtNwE3ycnaz10aMuKzK3H9Eo+yzpFG8HoiX3J3VlSL3TK6AJwHtxKgJkvIfdIg2gqVp/nt
faVVtSyvqdLa0OonjCG/De2IksVewlINdA3DFOmnbroG4xWfKcOsMcUROn6lP4llwiWBICbZidQ7
hU4llD6cv3plT4ky9MeQznWz3O1yGeUizih0jsEYEwX1ac5ifUeLXxRA/ZxLpFOOHwAVHhw+mec+
VXIf0HoFqGD7Efc/mNZnxCAWB44pP6rKptTzHx5ZTIVhZBc391OEekrpMSStIgepKs78NVbRLSx1
vQQuk1BBEeiC4ergrOVCPnMNchSEyILiIMP58hxn7ysZrx4pMEJuNNrprtrSJMJKR2GH+tOE0kqa
jxwY4fzYoScqKFXCRk+bcK62yBr6M+UYqP0iRRZ36zSmZA1dUWcrVzB6jG5lC15lgfH/q/F6D79m
+epkiLSR3Nol3GqYFwsio/pFBfVl+eeI6/fjn2yka49IbIp5AAsUOlT/7/h/uIEizZsfi8bFZp4a
8zRzaFTkTwtwrqIT55VD7g6X1cKCnXfAvWsE78H039BDB48xOWiI0Wvu//z+y8bumTs4gOklc4/C
RwxRcCxWyxVqGetpiIkOPLo41bMyM5eSGXFixdsMayJijTr1TGHHoUALM6HFdkWjL4WQAv14P7qW
rF4CtduKBy41BCcLn8vFlNdkliwIvuWLG7sTiK4asYGoe7bOd3NlngpvIAsQ8Ou/fKPHlNmEoYR3
QQJ7ACohCQqsDa/JMspKDHBghdRVyVw0QWivPAOGDLZe9/9PuYh3e0Y7jRFqVpkVzsl0QAHGdV04
qrf1HuSCgBnOqRMK8Umg73wolpeTJQJTURdTTI7O/OWzZQ9T5ipnZP3h4QPtT2i+21k+flQVMz5k
PlbAVDosoiSo/YPYUbLuEoUdRM0oZ/e/PbhKPVMk9SfWGCmDkhOOJTw8Xgh5tpvqUerLYNEQZoEZ
wk2fCnTJ3aJzQQQNM4tIAJR+m2NU03TdCaH88FMZioTVpPw+hEHr7rjoyxRkpwGo7uKSh04ZnDVC
gOfBXGKjk1TdrbEzkWBQgQNFbRj8xfI1p0mvw/7AFtU/O6fHdu6HOy7iTDoUKVbJIaY1SLu+AH/9
ysC+9RySKM6sxCUnuN3NIH7/NseMg0ABD3RKCvmsgfjbjrPI5I1zEbcfyyT+9zFMhZ5o8mRjDYMJ
3ThUWPFJ6BuFJwF8xx5mnupfy9NHrx+nGvrXDtUgUMT/Y32g05CBXc/DPLnu2vp2Sl0lnIE886Po
1GwFd+vXgdTiGX2tIFQg3qDv5HpV5oM8iGCk7/43eES0L8MspU9ZTchaMpFGKdr0VK+j2V50/XoG
RDG0fpAYmcpEHhdBs0wQkFWgbtVDTBCFqNDmli/YEk3a5uxs1r6QRMAaHoIQEo5SgrbZIw9L0j64
MJyQrgE9z7fLnMo7M9gAPebeUri+Kg/rpuBF8gOC6sVxvsMcWLrEm3YamlvohkCf7HZg6J2un0DF
cpidiYUfi30fpIMLPE7vVNUKC2akXS8bQzjHYjwZrIsmI+4pvYIPq9M5ns01Z7/Q3kdsb+G3Mniq
2Kija1DomosARnExd1KuHMS8zMamAGcBGb8LctnqF8T6mIGD1QQyL9Xdz9HbDrnbX7V7mVgii8VD
ehPSeNiZhZu7RJnofDLc/ztBBcQoW4KEDlRMh5EqXthBHBrEw53wMblWkN/uoSna8igBYgueKWbG
tzttuGmardWf3RGrdkA9w8KZGzuSWMUEiJTsp9VdTV5TIzER3gm25gd1GfvPjmWtSUn85jyzbJ24
w2zR4VhGf1ToAVuJGgWOwbJnQvw5RH3cAYsor5f675aX/h3AF+Sb8/G6HizBsu8UbIR60cgbf2eX
+jqovO1THYWo8nywbwGrB2jwiNR24+IXYeOXoM+Szj/uZvrElxKPCMcftvnBkKp832iYWPGxdNvn
uefto2gGjVnImaJEZAeJ8ncbChBHlLc2ujldVsDjMbyI3pi6bmIQWOX9KLS2+XjDHiKf6mKLRTfz
AJJq/tvWZeuXiAJl4+7yq5Kwn8ftObhkh1hjjGHKAkjSA1nFf7RlnhCJHEP60YgYPBGPGwHd2NVa
+l6o1de5BtCYW8N9hQ7A/NwpQ2rQNg+u+k3UpwagwOyqsU2aFNeLjq84cqtdjSdOFB/Ce6yQekF3
UdqPaDcLHPLFMf+kGumtN3HpWhB0zygiIk0Wg+3oxXEz+nUQZE9O1t2rfzIs1fO4IYvPn3+5HZQN
sn5e0F08z1zXUSZjLbzq46VgJAeT0dvwEthJ14Y0EU3nNxg4R1AT4hyxbBbvvLHif6qkPvTCz9nE
9YM5Vi2P076Gmb2vLZ7qRpWihbch86wKL8XpxFIO+DXJKIYV5GoGp6H1EN8Wy1XZ2ctD4LtkYDmE
A6pvDbTBQ187GUcnLTB0AOC9fV4BeMc472oFKpf++ymaKPmBLB/EzGX3V/KlIfy7gr9S5sX6mMQF
koUQKkuHby3/Xq79Tj2Kj86VjSBH3me+yGo1l5LUuBhRMP6ZOutK2AREI9LYO2zatif4eWalQZe/
A9baMa1etinHhRqNLtwZA0jJ7kNKy/e1lhnaJeNko6KEzO4Fv8qcRVXKWXqeWvEJHN3T7BGNUF9T
rTx4sZddkgfeISYKp2iKWHpHxNftnMTlAjeF/v095QKMT953nO4foe9KFreAZarbBB/hbsMUsZfm
GDFzywf69cDNrkHpO++z2+Cs3onZxc4hRgKyZXFQQwoaALMwFcY6OIuZlmwx/avqVMSXiPteF5Ll
S1nLu9GpVq9F1R/L902LmaGNafuZja4OP+EscHqlT3BqTN7UCoOiiEtVJCfbeKnLPoZ23rI8gfAy
HnDBzhKo6VXzvuSvB8TExYD6n4dWk0uHboKFt4JP3PmUvvS3iXNQteg5nI2RaLQUJWqqIUtbVeTI
EmQ3NAH1UlIDkOqqVoSbpyj3dtmvQtAzD4TsWsSFJFW0FUOe8zTK4ndYt8Yl0KCwuEWqhU3ZXsXQ
ou3HDoprPHHaumdHKAzpLTZ03e3ZWsNYvqSmqswRMi22+Hgo1AXG36D0DbJ5flA4VxTqdOwSz5ys
A2eBCyENt1VCBtcT4G5lrqh+zSoP9Uvaa1ID2qQfSgO/pUCB6sPVkxrULftmruX1o6tWt1AXldQl
YguP+lH2Xk3hZGzf3PbWz8vgg7+IXY44aUDAOoL2LArnJNiufoW9EJHO3PQg4vgGLLv3NN1gS0Sk
0tNRIip9PS+01K46i1YGbj01y6hwM8tstlc3kT+nTpAarxCp0rI8GY+5BK4JCfqh9yoJC/mB80j8
Or3Uzwzdsy9OmflDI7OHA1GZ6mkS8GRgtMCX86CI0LmrxwNQDrE9Q68xfaiqKE7PHwT5Mg2X+TIi
zY1Nk0qBsfmu+ToU8VZ+jpq3zx8KEkvSzv5gpg3xlVwc27qDOa9buIHovNVhSrfV1Gy2e/uPZa8A
z3/ckezBX8jrCBN2dlNlfZXe8dBf0UDQusvGvAan6KqBRMFn0xQZjdITKLRk/UwdcS97chV2FHQ3
Jsqfy4ZSQTkQhJ05MTbuNaftCv5S357P4YIWJjqXGA2WD1kfzEeyFAyBT/IJO81+zLo4g7dGKaBp
Whlf+4sCAidqoKssdwW3E3XKeKEhsQ+MTuZdhCHRdtYuzVCsjAciZWnqfet1iT/RgG0R92LS7wQi
tQ5mVJ9mx8YUV5qSigYZLmW91WECeteg+7q+Ddh31sOhs+z6Iu+lFbJFP8V3o8qKcTJ8iEchJeBt
RW4a3kK/Fpz90xcfUDaXBxV3U0V52FLYiuRkSWqPn4O/0YY8ARr27LpY+ryCHoxnH+IeI3ArrJa0
3CrMxk0L7EoUkE8DVEPJH1GL5Aj2XLQsqAIpJi8XrDNwqfeDHIy0ngH5NQcj86Sc2/+MwIhV3385
hoBTSSLWy6j5SsvYAsWOKlXPACBlqs8nmKku7EEcanSLSl2Ggedr3foiEolvQdb7igKL1dBaJzt8
3IVS+Hj7vhCnAJDaliSRUEpkAxiTlH7yTYs7mGcSrR4oKxOS7WpLrMB+IYnWxLOvaiaCeN7YetHH
ffnuQwkUlV5NNhbskPVVfI/HeZKz30yLR4uCNEf1FB5Z8Q+IlLi0wIAiDSloDGZFlVlAIEfl65nP
qElUHx7REWSJdXe51htZup0+vhQ5a0iAyASYm0Mw1a9AOrQJ3ys2Py6TB8IGXK3EsursBFZZ1xK9
NJ9ILBev/Gvx6tU52c6uUscfAl3efUGfWNydiI0B/NrBXFXHXLIA7RU/8iO3Zy/9BtD2mv6R7esY
75QUDVECTQR1ocaaUP4qVbhTUkk/w7XKJDVRfsYeODP+aZFQbN1xLh0FBY29WCxJ9/kOa1WHDnYf
kYnn0VlCXhyyN1XEoTlJy5JUAgeC2hKSCOJso3xymT8sj+nlCHIdz7UEspnOPpH08pMdJVFifA6F
zvDmVMarRsGGWpZGrQoE06YVdpQdF8ruDJ1ShCYbJZ2oGwezt+6Ki0iAk1NM6LhPKgjGU3afKCaQ
pclA6vIc05R083Bi1Sy5xzmcTvzkwnpWQlhjddi2MqOt+YrECNoZp2pSN+yAgOw03WBCmpwFaJll
PFLaV482HJKk8ApbzOnOmV5RDQNPijcqSHaCybFJ5znNAhfwd+UomMuS5b8fV00daN2SgYmasEC3
TWwL/tJ8LzbEJo+Uxi2HmaHhbsh2W7icTQ8ECe0ou7E62Sgz5sJZyaMxHEabKieBg0K0z4OcTgQx
rvtlCtc0HznuuQ+UtZKOhoq1Db7Xtl0ddDRKwcYiwjsGlMfl7osHiBvPy9PwEHy9jBgvJ5UJi63B
FJLQTeImwx7lKo8Z9P5Sz0eNkf/fK7ku9W7n8zy5j5c0KpFQ2p8Lg7Nij/+XKN/RAPVuZpiOm/fV
b/oHThVlPV/Hw61Id1jTNmqBnwa8Jhccw8Vz6cUPfTzFoFOnAF7taBVDfKtkcVK3ogWUCePAn9W5
ob8UgOjbyScnqNE2eTbCnKZxKZ4yqg9fQGXbJHNuFpafjNmVOb23vCuymQR3U2PgzXhdM3QIBn9U
1unqvtgRFqpQbYpUAVsoIBJHaqxoioAC8PFI5NAcm5BueGr8iq84e8Ode50FI9SEZAtII5QleEZ9
ZN2i+AOv+p2IXURPwD86qXdf0pE8eblYj1OZnB9VpmbgGmhudeNXadQo+ma8j+hk2qXTg/QXcgr6
5M79pb3AcsLHF/sOZszH+Er+e7HghjDc+vK0Mb9Cq8BkHQCR7HrngbisK8TY70OECAIztdohC64y
vYrHEBcboSZOjc9Aq9pik43qIxfZ4kGx9EhkrzPMmlT4bfC+KtsPMygXRdw8JWXK79OQVrn1Dmjd
dqj07gczBBZh/ELB9Svvd+oLGceLDh02w0hjxvvxsD4Dh1BOhTKlzNGx/96F8JIuqm685mnj5K1E
8VT1iHfSsTvmnVzUnnVm6wM9891r2pBt2LgEl0xKyJ+KaIE12sADBKY5aXg476WZPFKrvlNnvSk2
h2jgtMmWfNqIcWkXI9B1CKwYwRBOtr6Exvu0XfVpHs6wQkRoZyDJ3jK1+U4xGhwHRKURPFp/6TIa
mcCAgfN1y6EZPFMX6W1r9s8LAv3RXwkwRnXHMTtKHmRrGq2dC7x0idxWPK6Qp2LDumqVcqQU9US+
E/phU9aOOHHxlggeizIkpk+5bVRr38bt/0U00dWjR+634hybn/swpSACczx4NKtXl4EXmpSAwVBM
KgZ6sv22H7/R1uQ/lpwLt9zEWZFCqhFrX2Mjj1AB2mrpqonpRGm4wj+Gr098796SugYx6iPtitrk
Uem6nIo9oDXtw/manEDB1xJQkVx15ztJvR8t0T2inL3xPbfLtMsQ7/yjrAPJ5SEV9NRWxA8KSWPv
k6jvTGt/EIjhf5o59TGg5CS/+S7gEEFfxqqAqx6SaOnvTv1H+hVX2gh7AXyYPSNS7tsaUCTxmyPe
HdkRez6Vc1s5B4XREU5yYwErbk8A2qBZKN8RtBpJNZUh6nL37GzknrGRAQSVcoWkRoylVXNebCsH
hRDXYwcCcp821k8N9LGkhrtsBPeYBK+2Tej0BLaDRR8QWNIWgXx/GYKfTznWJYEg98I2NrY7Q8cV
HHXbs5yGjwi7KaSvEEDt0T7OAfwHhdjpa6bTYDEUIdCOrHt4yuQP0VlLL0XCu/Jgm79EqV9z3saG
SygLMv4wJPrpLgmy9mtABjIndDV/WhAcRA4NLZFurF8oXA8U9A7OrkmPeboPyY47HnSt0+hnFNL7
o8Wmffg/4bSL4POjNLKnSIM7oxN3fhZaFWc6dy7Iy87L3wJTay1KR41NTvPANWKj915RUEFF373/
eWSLVzGfCBq0wNf3IsRHf/vxtbHu1HSKiyQJljSPAVZ4/GWkeOpshUhOSjNpxLXQxDngwLc4AOJX
kGW9LeeroyrCKEDxnrMWJUeMK0Xpi7Vuez+WqF5dIB3C/C9voxJABsBebOV1onYqwE1n3jwSbP1C
pbbhl06prdkEGGG7mlyLQxMxl9k5h41ALMc5Bf9zsZYh1BP2tBKbxc0//Oe3I0sOMhoxebkFtbbK
UWqOPUWzqq0VeAMDmW1YKnmBYmNwxBAMNuV7JOnMrq1BwYQhCVcUb/VyUiSjOS22sJgcJmmnSnwu
+PJBI5oBcC96IlT0+M6iFxifu2yExOsePUTT3xY4O4LjmSk97tnZIqSgj7EPl+2C6CMpAuUUakBp
JXWIJHtF3FKXj87L+Fz6hyjPw2iU0Auizou99uzIWrzvhlGUkOmNwYnrmUKumYkUGc2cdYOs40Y3
o0+jhhj1wixjSV4iaXhxP5UGFLjGMWoLwU46PkmOi2qtJNdsIcD5Vhy6l0kqFLK99i5tqX4FYLKU
gAqztEMW2Q+IbwwL1YyVptQphQQncXoRAAaTjWdaTr9kvVHkhiVT3BcnsFfh1IlDq+hfxre0gc0i
d6OWWueCkKPF74cKygd3tRvk9LyVrRJELnRpK6Zz5kpJ35m2zyuvbHfXdz8kkXxiDJCNJSaqkdpK
jEKgtzd09Hx5rF8XRBFrSj9T050ile8Gr+ZE9R/DMcBX+wB8t82X5hOzerqh0d+3q6QyHDkj1N+k
5fTKSrd6EVlMKiWSNv7YUIjmD4mNEVRPGZ5Bqxl8nHOcBIBeOmcY4d+RxMUlJjPClep1tV0AEc3C
RnHEafc7lxC2rtAvIohuF0yI4T+XNyBl4IpdOM7RAsu+XnMjVMdknz+x0c9m/OQOsG3IBRr+JIB2
/Du65bjrqpAEBIPub59mTsLmpd2dFdB8C4JuRLQxlzI/iROIkb3pk7ji8BtIWldpQQCC0E/iW34C
iKSG0qaTpfVdpRsLpDjxTybA71wRDFN2LYHnEOzDpMo/UUrFgWkf7UGb0s5ZcYOY2WjKiS0/EHkF
gD3LnAlXQ5G/2yrp8SSuIOeM/dxx8+pRUjxYfkcKbQGWn1NYy1RNAKRqb9Vm2pARtFbkhPvX0V7c
e1J2Vo/G+f33N/qTAyG0+8wjxRZR9AS2QhdlUxuPXtfChYZ9cRPolycOVjbsxXwDqw8DAtoiPoko
lz8uxXmT6AHFP4l+No9Ka3mCB8nLcS97+4dghQjuPwEHbhx69b6Szpt4JnL8y34CaNckcwFYbpNW
QQrDWbjV5xIt+64/T+e4GrRaPbrffRgJMYWtXdTaksN9BStqxYYHAcVbDNnZJRF0quU6akABZ/eF
r5OsZ4g2CD925KgIru940my6/MRltufmVgpP6zykSxVSmAF5neP3zPAc1ECqfOcQN0I6f2C43X9H
Jx61MR08nnpPkuY1THz6O8Pjwb3zHp+ONUoXbvV4XBO2T7euYEI1UjORzXct5ULmWZjs4dizmkKx
nDOD7HmDlSeWicmPiWrWfUHkfgO3OP+AydSdfnrIEo9TVh7RkZqQIBgGaNzEnoSFNqKJ1N+UBauo
VsZiA+8FtiMAsglBj3RfVl+dXNXHSriKlF7mmHDxtFZSNb6kgz4piRZg8uAGjFqWyIiTPxhZrUvJ
AgA/PowcS/a0tsCM+cYPR44yIzAthFasyzcTOBtnVIb6DSYEvC1nyV8LnUw/3cN0Gsm/rGYAJHuS
FTokhHiKZXXARayuj/RifMY96jkVnohgPSo4ZqOk9BrOL900/Ulgx91tajO2WkGjo6RGHiq0fqNf
1MMM4/8KMdc5SJmypCNtA+oVJjpQUQOnzGsX19/TA0k6xZlRGlqEAzKz6AOSLSVbiBPXSQ6W9yCr
KPbJyIE5n7sBr1HYlMVDxVF1vTJsDoi39ldoT26m1Qp6Y1gbg6KXQuo67zhHc+N7sm0YXAvP6RKO
zSKuKQ2oXdt4tKVLB+nJBlTL6VaVckcfWtssnInLUTUVyf7rha9SKN1woTPY7KFEsUXh5qDK4ZLi
ZCQNGAjUga1xmtBaeQXcyy5JWHEo+3V0J5V2P5AHm4k+Mhp7IW+4WHuUUJHIgrSixcTVAMrB183D
dZbKdXINjIGaVRDB1XwN8GHOyJ0Wo795Sdl7TkqIoo+jnfFNynKgh9Jxk8aV72jefZ/pYEksgGWh
UO4S8uj95J0LdjQ/NHNramQ+FArC+aZciTphacM34BFRGAtOSx81ZEdtlcY0gOFCuqRcVp/NOapp
N6v0dHCzp4DQjtkk8Us5FgR374RmGBN+Dt/V5gC9dKPpfAk3Ju1QLFtUFklwAbj5Obh4WHnE5W3e
jtKuEKA8c5yKqJ8XDY3/xn2hAekTiP6v45iO5/RE1FFrdCFiMMc/WFVrGMHXC55E2GbuNdB+wbmG
8r5cclEdu1Q4N3AO7Xe4JhzSGxm976Xq9TXZPE8rbimDE064Um6agXGGF7ucGGsUR6/0CWzXN9Sl
bMihqef1BifWPYNtW2vrApiclCmC61eto4DpfZiuOKFvLVXBzzhVZcjoiU7G12Xr/OpqqoMM5yrC
xS2rHhWvWHmEd9ydF0nErWi7gF5rp4kYrhcBstky9NZ44FQjlE5TsJ5BmnESqVYun5+C8B90GxYK
5eupDIwTjVBVBBKlIKCKWEbzM4qch3tNAV4mafcy4eCRLDNIX/dw3AMoFZT0MpnIigmviVWWY1sx
wCEF7D47P06j+W2XzeCkNgU8ljogltax73J4cml7ScVNKcGjuTjSA5OOrqoAbKfdRssTdCFXDDeH
NZYoCiZSAAF7D0mOqRtNs907335gYo5NG4XkxT+ZZNqelU6jbqezP9i0bcz8/tUZRTa+tJ+TZHkp
4BzIDDvSSm7WWupYSShBzm3XG1C6tjo4AOm4xreWUSQM232r1x6ovI/teMOFhjHKHM/eXJIAk+4j
o4aVz+OA+MOfX7tC2G7e15unscR6RA8/nBYZtyA1eNFiHfI1CBeCHW6Dr6rLJunTofwt/+1wSciH
FZrbXCgKxsuSM1pxEI786LUe1c3SdCub2FgUnCvn+2/sbl86cByUBkrJjyrCJuiaWD9hVZ14ngE/
SFnH6LnxGNqCJejK/fOi9QpD/qFH13g2vQE2pd/Ex/f0avTRrd9ACshDdQjSG0gZCX3pLMfzrK27
Ntyvu493/HPk1gKLVdhSogUdZvR5St52l8UmdR+JrcTNY0arOUUPVdqzxXu8ZiT9lt44OdPoM7UF
MKBVdHYJcPenIYmKaaQRL8YFqQ20xmc8x0cdI9w4pl7+6B0JcvJMOdOM9U6hELSLDq5A0dBklFnm
szVUoJjqYMeEu9oZwjZXjmwXfVSKqPoBXTUeTwRrBz+wXxq6cFiVY7ajtq6yEDyGJOjEkteSrKNr
P/A7g923KOc1VdF37j73Ij5tF+dZgE/92XYZ/hyuMhQ35OvyTLmIntyORK1H+bJLsLLvIyuimj+p
Ac9jjZHkpWUwWy4U1HVm2Q70Ne5FiTB2B8FvwjJIvs9y4Ct+aGpTbPoq9PJiKE5Z+nCEvT0ZlDr7
5Z7Ebrx6JwR0AoKu0jLd1NO2E9d17iMCGZbwjm6AOdQnLZ2GErBQ081Q/UmPH/YYUldcczQxgz0R
5k1qs6z0980tSybCWmB6m5cudedgBk+/ki5uUN/Ht6SYZobWNJhG3fp1862Eu8/CYWHu9e7pBNYN
XYjKVH1Oy9NA4XE8xkrEepFZCGfuFQDl5F7a4CHvzF+tURWsPI0fiI07hQaT0LIqjwm+CLHaNcfd
Qzitlxk8njh+x3Tq7l6STYwmDGnatnFgpGDRTQD2703XiKtUWUEqOz2n+vx24LeXM6UL3sMkQx7p
eHGeCzLBtPJQ2KsB3L2geZYR9JSHoMqE4bcnLq5tmbxaMeWgy8g6OSvz9ccsq0EuW+Sm1e7biTOD
bbBFFkJnTcSaSrjQhXFga4gUIFMmS5r907Bmzmbv5h8QuuAYiiZfMBhGcdV58/wScNY84jvgk8VK
amVGNnPFppIv3KfB8eOHzPLAmGVD8xTWIxEbeKTK+m0XrW8ZkjibTX6BVcZCWVL0zlWMY0RIarON
OFyTmqYkJtrUIDW8J76/d5M+adyeEeFLPkrmsRzK4dNHUp4PyIRApGmTrawqHvc6VrlZu4e/YOes
sy+mnNZJ2XFhDF2XXqQKHuprvvxwVd3WBxT9328ZfBUCxrGFz+arwACZdqTpWh31f3xOPfYgdnYL
if8eOvAXaQWpnjPnswSncdMl9OVEnAbDNLdag3bwhfVNdgyZ75B5Qz98O6j2AG6iJlvUK3EYjLEQ
A/7TWCn8oLkPqaAVsmJm/IRFtuakg8yF4XtsTj+05DBWu0hO5qCz4dTjwpWx7/xxKuaQMvIb5KmF
7s22y0n4uNMPJIlwIKYct52c2mrpoKH5PI6CPxe1+pU58dorDUeF+cgVQ9rvDpmfLolWCwZZUo9e
1K0rTytBfrdSWtW53JhUMjoZcvnJz/KFh+UoXvZ3ZFeEv/cRLLB8w2BQww6DZZyB7FAppcsmto32
LoWBoI3fk0ZpcDwYqO6A4ZDCmOHRzT69vxanxbi+uXayFJVvo3GEjwicbXFFcVm8Af/kJSxaErDU
O7drdUlODjYnQW/oeGYW9LoH/X8/EcM/sbVrymfsNxR24cWNbahsE4Lazvf16l8vBx9xzErZUOi7
IhD0nbu2PViKRaCgj4iDRahNd+mjESX+1zpFwJbOY996/tVNIoIXXc8UakOES2HnbJ8c2bXgnr7P
35CN5h/TIWnGMiQBuEcmvcbKJc2S0+cx/uTAN/X4CCnCqmGj1rnXLTbui/Xdx3sJV2V0rcv2H6kO
nST4foJiN8X+4gOJJdQYLxQzgpUCAZpOFwyIFZ9hYhl8BSMjFdt6o7k4cXbqWdshlKtRT8XsUU1H
m8Yrv+swYaPtftWfG7t6pxm2oCqkvgVNlYLfTG4GX1heKS4VFh7AezCpQnQe4a63KZ4kl7oYfqQ+
QCC+NKmhau7Zgy0Emlv+RAwTGLSfPWJEe/nXlGITMSaSrJtVgPzFvNRR9J1HL/oZasjL4FOntdod
Y/SoUhlfme9W8FUMUkH7oruWZtPZMEPFFvbGV5G8lfrtiEdyXBte7fHtwCAHentKyKvs0Asj6iSx
zQsoyHlvVoHZfdq4rFVC0XRna6icuEHobhvM5ylVTjjX1tgNdmS1dmP2GQxtVKVWALVK0Sea2iaf
Xo/BsaPVd2NzIA34EcqwcU7mVoGZlCMMB1iaYGvtCPT7VivqZplFCObOWLyL+nTMPJc8DILMGDvL
MuAUA/dvYsF8nYfT6DqggP8rdEzuLcRkhA8DHJ471NfH09WMkPVgiWDOreMc0A/4OlASx6CfsgHy
PV+gnrP6woAEgHFpLOA/I8Uh3ew1g9zLCk3I5GW6QvRCwj7w+Fegb5gKoUCw9NYoz7mgJgonWO4+
1pcICTtTu4ASpa4O+tQLOtiRC8bF7JGHgpa7hDMSi8725HrZVoPc6qhgtrFrDNJjPVFbkC4DRA12
Cql7nZgkmiRIeWvQKQcuUr1o0658Hn9s5e8PtjE244ior5lu2prrSbZiOmjcXg7GSCrL1oKmri6H
0aLTgA4iydLHRgXGp0fWWiLzcn8yhge25dho7SD7LefksWfKasv0hCMTZy/PV4gvB5fLEtNGyn4r
7TMOoJYYsBj3b+o/xriuV57dNF33/13c6MGZEEURO8sWU7rjjeNpwbLsteEwjB17QJI5pwKcAOL/
4vv0m8/XM5P2OH/dCpkuaACTdw03r0jZsjWbVsRGQvo4WOGBidfIwl5Fl09mWFtD5/ZkQRoNmGct
VsO9UGnaaSrskQlWbYZ3gq3zz9rcoOGK8fVoiTJ0uKUeB1Np++eZMcZc7Bl+6JbvaDHuIJKizQBF
XVG0hJvDCDllA/PvKiOwAkC9ph3mNONHuv/F06JCuHKf2auH0SX3tn6dTAW/oIVRXYdQIW3mlft/
2P9oLzatW++eQyccH115kJm8mfjKmgCc8ISR4IG3VjKyJZeoQx7oVdgfPSOvhLVliC+97uH0TQ6Z
bL2hbKO7Lw9+TOn8mACbOkdJe8pkaAKrsvrsb8t3IrKY2upb448kWMkN4FNOHeGYt1/UCI4WcY22
32HAPdgMt7ng1PDyz3VfkoF1+2QnuhOveITcIRGuMiC53EPFFOh0D5NjzdOqox6e1PFZb9KRQFWB
dlpxn6MujyOOHzBXJnZEkI3+7RPW7Jtxjk7sAOL4qjtJAiP/DmB+nhu4omMnDRBJNZX6hcVtFSxO
ccJV1vuv58gdRcxAHDHUbisJo7wKIFTJTeGE0DzhqhlXcdQ7RYyUi3qjaGrJKvFepRwpN3mkBWhl
ZoeFcVZ4SEjiAmmCZwk4LbnIBoulNFt8Lf1NQiwkRqZbAMchqJV91ZrFCq1/erzmAGx8NRnpVIWx
0PNOAvUopwZz3JQKPtYZ3U1Siwax6Qu/UqPtgM1UIZLkguvOfrMInBrK3Z7SCLDBqoHEFy6eB7qM
Xb6wFVrfa89myjxrDskZ6QD0KCygg4TyM0R9xjBxU6RLTYgeh1DXmTr2Y7pA7LtIiRf/UcyNpkbZ
onXEuLCrXBC8SRDSEJlchgYC985QyrMOrjPJhlRh5nl+gQ4z11LX2NDVSjJ4KKuZMlrSjcQb4xYw
QeH9UOfxY+7D1N3cGZyGmspfBxvOmoKcC6sDOpjsnIJg5pHivuG2BJs/65//R3EkapWBOO9M+hTi
2M1V2ryCg6OG1pvmWOfUo7LqEM1QcmjM+1g27pz/mF1hhweQbd+OTfsyH9tw9VayVyJhWtbIQ4bc
nmCz8QZjXM3CTa88s295si0OnS1zOmDq+Zg4/lqvdBxhT+BbBoLeE8Ce9L4iZtDuAHCNWQr+6u7n
pue1WDfnZqS0aYFHFojoTlUoQcI27jROHPyKfDL3uN4BlGBT6nwr6DbvgjsMSfni9SY0OHZafrpT
PZqur9dpX5dSBeZXUR+Pp0auBltpbLWgV19T/tEu7wCRW99hRvSjkuiR2tYjR22mejNR2szF5hjL
f1pFTu6L5fw/qiJ4v9vkBlPyuo730MfL9oQ1dwpGgyzg0eNF4RPEyXo1c4cRJlDJYt5bpnfGvO/2
9e8qeNxm+KWcvpqNPBxxDJzXoXAZZlSxJpudKZrvjNPIEVwlIVIYTR8ewaZn7dc7TLvr3H+/MXZD
PaknDtjSxs9q9beXBY4kKrojeCDKdxfem4///qvgYq6EciBIEMxByg6J1l/p9z4+yEgD8j3tYxxd
8S86c4LVYuF3TrKW3eUxt+7J7OkH7Dmm7aB7+PvfB7DYPhbVmLitP2ZgU7rLF4f6ryeYsrvdCbin
5UjVOlJGh/fEWuqhUcQSDGT2rfazAc10mrd7s5wtiHoy11pYgsvYp0NXDkzBUkOWKvCqtIvqHorp
Ui6zRC+0Aui6sO9TIFcanoGrUOrwkE9QO4wFEGEA215eKlQMAT77JsDs7Z2Jxm5MKTHuBaIywO+b
YHnIKV4Fo5f5A8GL68fJYUgTo4O2auCwP64JbCva8hF81zGJJgVhGPsNtnc3rPKJ6IKkGgydg+2Q
9A33Hr3MY9Uy7vXfPoNzpQrs2oKX1El9HNNDmH2fDLNf4+O5ZtYOczmpLWJqNcgb7nESZBcX0ztu
aP2zzueP9RZexF/HVtYu7OaT4PxB+lqT7XuGZN73jVbJHZuykUSr1uUvr7wSYoXWDTrfyHgJ4ZzT
OZ6owjKaC6l7HLauUj/SUr1iPrFxtkihokVdcqH/USXJIlL3mE2yVePYfzZlgyRBhlsFO3WhemZa
i3PkFzJhWqEgrYlssCregj1j5334Pg3AVdMwoKH0aY9i4MaDqasZ/ozjGLHoQIA8BdiT7coofw5P
X935gq9b0iuwgBt3OwWyFtbEZeC4Ocg55HbgB9xauaAVImCHOQH0z2HecO1wZMuRAr/mDGgznNGN
nW6OGE2ahPj0ToLQX/pVSfaVAm21uipEIdzoUaNFm5zI2/xemuVw5/L+SiAVIO63OnjIuWz4B+/P
9/ogkQ1mzbb63SapjlG+IcId37i3ev9dll00s58zp9YmssKMXZu5JcSFSKfQWV0SonjJiC42SFSu
62jMr0nORxqURjZiKhok8/u+PKX/r6uqZ91p9vTai+ym2EF1FxbBIt757mUT6HMDi38uCSvubtd6
4ojqQkY8eEbeUA3U7gHgh1PPgbLAz4wFbfgY4SLxpqGE6QlB6Qup+O9jLCHy2kCopvMnwHkCHMlH
04fe/n7x03JVLlAGlPHlk7DPLH5uPJ1iAei/KZtbrIPp7qslVYm3pOXf/X8vf5Litq+p+eRSw2KH
GoCv1HFdXuXQq1uSsoJenbw3pNn6TWuolN7B1lOPoIqp7WkB94MdfCc9LUCHoAGqSwMsa/VkTsPj
7vwnoM1QBOjJWOtct2g/Vicvge0J9LLM7Oe+4vYn7Abyd8JXRVbifmAXldl8zJW0KDVHOY98aHHW
X0EEyHTa5dpG69nWIdZ83PZzAkssacay9nKkMTxfGQoJkmzqPHhHwqgUs5JjUDNf02CgT0l8lY5z
kj32hDsS8hHSuJrpGR1s5aXl7NAxY1M4CqDg86a1jUJmT6fCDNJASN4vnfQUIZJhySeS9f0xDTuD
mHMIc4umLwicP4E2flgkuek5daXSyCrx3qylwOoPJj5xCqy4sSwslG7NEUK4jvTJfH6qwqejmErP
IXDo/4dAacNQATmH11wDmJT+z+EE8YbsVQjnooyKjiKcdhf6WekPM0FOZNjhCscVZMNGiZLhZD2h
wyh2IpVjYCdfVc5wj4h8YUrGWFcFpApraQNO/oeleHhTiUAmds/yHlp9XB8BhJCkL8MdSMbqrGqq
3yGdQpJ88qHiq+gsOTjZFy9Cx4ws5DEAmDZYN8LDbfrm/O6QJ+mwEXG8LkOgQmaaeid73omTMfQS
hShKI2J0To6mzwwuuWInNEc43+ckiSPl1jBB8MOwRpI0wN6g5m7M/2aSFMCkJw1n7tRhSbR33oGq
Vbuiz1U24eGWs1ZxUZwkIA6WrufgOqg4SxiqfbistHUBZW6aSdZ3KGyLZuPZSBUy1iwhYTrTP7XZ
fFqh4wj8o5ajN3NbRd7nVsCnCJSeHJP01AWPONZht/JiOtpnwjPA/SdYosLUJBFY/vZkWYbqGVxz
GZjAtVFZnngI8iIZI/ypcMzSnw1NVa0pJD1ydmevZipvMe99WiZqh7ZHdb9wuDRdKfbOiZcXwyoj
k8gkrpcIwVkrDj+1++XeNzDoVzLJCV6hbGemNVaRqDjhx6+AGVkkFcZVFjj7ZgtZOc/mHHgXZxqI
9a+JeqWjUlscBHT1xLGIH6HXoF32eBCASoq1N9BZTHIQnnfouSEydkYxtZbLCL2zNP3v+vEzr6DE
uPZJOgNxTnl68L9RAuu+HkQ3nWxNT1nS9sx5Q7QI2p2YNJhN8CrOfky5UTgFt0L/+l1F9EuUpyzs
FgATOp6BUMSIUwsAa1DKTfKHd/ymf74Yt0PTZfLEYu5+7StS9UyVx5UmCRr/OCjCiXOkj0IcdPLu
N+9iFaVAVOYH5OW2pcwt16P8qnfYKtgEFAC6zSIWV+DzoQwwvRxCDFTtFBT+390AlDsBI/KmSDyl
zOUUYz8koNDucSBkbta8lmZquzRX0ejF105e23NL+i5mXgdrF0nfv8ZLucj43hzjVUXDIIXnJJ12
H3IWqPaYF8+yaSAzbKayE/32ZZFVavU0drukJAOsNwgaYTHTMvkXXwzqAsEmOiPwCgdp0Lpgjhir
ts9poOjxJtidQauNfqxKhmu7kgb/PXeqonXA5NoVYl/JiMzmEYJu/TJj5d/NBFVuILimffQLZtJm
Q34wyE2LynkYzmx/H9wB0j/kiQlJ5aBXajIVIUNpop8rlga8z9fVcJZHcX7DfCsFe/Hzj+ElSIuk
3DcE/4GFzujfDyzgdnl1J4oOnmv9yRAFGgDf4VErn+hld1qkCv7QwrhNk/Yt2GIdY3zs4wT0ZY89
wz6EA4VfJF5QjqauC5OGlFxeznBIuEU0w93Tn7l3PGWp4gNUZbaC6aAdKUPH9abD5887CxKas0M8
RDLIvBlWMsW3ItJoPvtXJ4SLph9RyDaGtDbthqKFLPV77YBigIU/NtY6Q+9Vlk0sOCKtD52KMvCy
epWyx70YKyvf8WO64TFTNuYZkSBpWANWc8sMZzgmHmJQojMQikGDkdQT3Nikn1Gn3b4BuXd1scbW
rEtW0Nxy9Hjf7uUWLbsGWwORA1g4suePj7DjoOMwHxmLL0mASXH4OELkb6Uh5icvryPUyQmhZ2oc
g+uq+GFbtY0vpeHLq8etPduAX+U0E+WQ6BXDS4a7u6WwCu2bp/3qjKduxSKAVtjysjS4RibLlTfp
FaCN81COraRNYAT9ylR/xbs7F875cuRNrbEELHseRpxLXJPfK4Ketsu5NEssBEWn8EC9GFtME9qG
exHVpcHXRPuJHjcDVeq10ZEa4G21z0KYI5iowRs+llzy4TlktNFipnXq/vHGXRlfdd6/fYLe102s
sYiIj908MdgjA1bzfQ6eARwkPb2yDtZopxI90LabTpUjh5Rkor1ljVsDZu8cMHA8acnp2eesXtEo
3AhVHKBf3HfGGD+pKP2c7Pt9Ao0Ws6Ndi4LX0hD3LWN5Jnd05G3bJk1tHvhQi8lEbVh6n0sfAl08
gBk5HTbgjyvcQQ+YXHI3EzAmwf4zQ7Ah9dgN6Qad9pQIUTvmJfEA7taqWOcxeJQC8Xwgh6rLtkRO
oNDj37wafiIkRqIH/x7apeKvVgP1Xq1PEopkPzgteNNgOUbul+ZZ9smYurQAIupE2tNZJxpgkdGn
OQdiMY60l9RMMRomsEFmxss/XK9zPt0+5qTMy4nIKrrUOmaONVFd+HY/vzqrY1NxDFJv2N/5G/sz
JwL3xGsTKGPEIsaqoZqR/n9ROg8N+nVitbm5DakDr74B7wTakMyY3tCLCb5pvMmKpV7YnCIHkNgx
Y1Vne5YzQM4/fD5SY0OOcggZCFH1X02AbM4+9nWIgrOMIAreyTGR6PUsOp9nLrxFLeh5Lk9ZYOKj
rlwro60R/zEMtSRAvMUvQLPa1ieKyVUU1iYlR9ClkhUySCnVUgameW7bVdyHXmuJF6GPdA7NsU9A
mCc4Q7jAksQQXi51OCZYSmHPbrwyoNEutNqy/HTlFeEPis4Il6EpRjPhmMd5FpJzaoOofPFf56ZR
HjzlDlbJtpw82jTFRk2ZgWFQIbNym41ejpSKgv0unpnKCJUHkNHqMctW0u/Klml0eEouaUOFG8LQ
x02P7TV5d/BA1FFG0IHPJi4lPGpz1Y+zQY8a5u4Vrzm79O2HsnONNDt0N1eTYKALXP/lFQ1AJq4/
2aWWSAI+bZsw2F6ktE3QoBQngsI3dTTej4ZfFSM02B/Ee0gWz1YVwSF4aCPKRrmi6hxjR5EdQJSH
PcO9vPhvnuy/A4YR4uCKLMFsRUVKN7VFRjLSEg==
`protect end_protected
