��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���/�����Cc��<Nb��.�x{�>��0����=�����=8RLG�h+OLزV����ݗ�@��&�K��4cbXu�6@A��?��I�=��O�s=���
�S�i\��D���d3�q	��9/�I�w`W?ދ�S"K7��5�,l��C���
@E=D��!
����荾Z�V�h��c,Dt��&�����]4w9K_9O�=l�uE�w����[R�\�zÚ�-J�$����åCj�[�
����T=���K���h�����,������#�z~��?�G���B�~֨1)��k��yq�$/ju�YA9��SX�{@��mWt������w�F��r���������O)�mC�&�����$��^_��|�����=������A���_"�s���50��-�ݡ��kVE~�cu��'Ah%�����v2ݲK:|�g���7/��=Q�u�~��qC���
qSa�a�n�m(�]�h-�FK�]�Z<��K�b�s��'�����C$Yכֿ��h|�[@lXJ�*Qm?�аR��(�v�vlr�j)ڦ��0p�s�bv��jy�-����(��N�vהS��Y�n)!��\|9��;#�o:�#��9|TWL��L2=�'���$ƫ���19�?�:H�A���T秧���,rJ$�p}�a�ڡ�rn#9���~�1e�[e���!������{�T�7���O�z�������쉎�<o�j��D�7��lS�ƃ���F�V�:¦?�,�:4I~P�o6����2
�ԫ�#��G롔�qH���'> x������>I�nN1.�yφ�V�ǹW�)��	�3���k��c�Rw�buRA�8����\��L+p����rw3v�FF��8��Y��8p��s3jL&���9>��y�(r�I)ռ��-�2j7�%�_�
z'H��߲�.���Z����k�4�}����N���Y|���9���
:��Z(�a�[j��5\@5u~�{xf�_+a�K� x�F�^����<'�A���!�qQ�zx�KWr]�mE�n9�
�"�ym�&�(�Q�
ȹc�@	��:�,�
w(dNd���0�L�V�3����@�Qfx=�aV�J��?��Nn�Z�
2.��g�	Ҟ��.�Զ��������a����x�*�ĵ\1��q�)8뼩\٪`\�		c�����#���<�j�;�s^�u���>�a#���.h+�H,!b�b�~q^�(�=�e�eQ�n���D5�nRL4@�/34���/��'(���To�����|!_JK�.jr���p�(�J~��c� �����5��׎F4!��f"�G��7�cQ)ܐAio~��z���几fE���C2�_2!,O���wpg�{w��vWb�bԈ�o��I��w(��m<=|u�l3x0��թ�˟zZ$B�]�AW��a�"�b��{��H�3c>���	�WQ��V���(�WucEi��
bo �p��ni`��mڨ��Pi����j�$��F�Y���"�R�})y� w���O�[:<#R����,jI����8sNN�?�hD?u��?#$��?��r��ڷ%%EU��v �s�vgA��i�Ǭ%�╃��������qk�i�o��3E39�M5���?+o�L�	��������>�[�R�z�+��XDw� \ݚ�X���R�^�Ϸ��Inl7��`g�>�U��֩�يޢt����=���q8Յ�eg��G<�=ca���A�C준��P���J��)��o�Ƙ2�(Lg�[7�k �]�7�	���ox��Mu���5���uG�~z�ǝ���_E)�����9��v����LY.���!6��Q����j:��� ����L�&�x��#�r�	��l^���/�\@EԒq�X�bNn������nb$eSFj7�YA�_��[	�9�������	6(��G�.�U���K�����=�{�!�B�մJb`H��i#�Z4���מQ��گ� O2�\�u�d��-��bT�]�xח�q
RB�e��?[�ٛ8 ^���PY� ��{0�R�	*�,nF�g���"g��g�X���d^"�,�+?uR�3|�u�6��T���8��i�� �� �B2�i�{=��DB���_��XN��rA����L�M�����xҧ^�s���,���+�����U�1$��W��V�PS�j���R�?��(��ݱ��i�}2��>��b���f��Pl�٤�qnuIr����V��?�|qK�gVC-�.`����~g��xK����\}f]���\(�G/���TO��8�'�	��}O4����{�XP�j�;V�G�0�������t�*��uF���n�@�{.�/S�5ֻ۶��4z}=R�~�[)�7+��iQNC�c�`�B<^���V$��֫Z����ex9�w���jE�K���f�i9���,���z��a��4��-�Z�`q�����G�O��z���x%J����ޅәd_�m��-Ha�Fu���S��!Ü��"�c~��%1�k�-lTX��N���z�x`�n[�A��.Y�O���f�fL��=4t��Bc^}�i�i?�� �G� �h��MUĸ�3X�Q[�I���8�&M����j`􂨵�.�m�ff�5Xe+��ZB�d�}-H�YF��%�{��xUJ�9�����|{ΐ����[��=��ƍ��wnHՇS>��q*�++�42��N�`�������l���Zf�SX���<�˰^fH?<��@��O��du��GAv��
����\��i�0�w�H�ӎ��N]�uR�$\�k�
����9�� ��eZ�[E�>
��ܼ�?��Z*�jaSJe���֖�VWY��%k0�r�6K�tق �ؕ�ǂ&�����^7�cF��7�O)xw{a�XA��ۉ�՘��u[�Ќ΂C}������|#_�gŪ��{-(	�G��>���-!K�o|��X�i�yeo�$� �dA������4�����_	E�4�2o�T�0d3��?o�tS� 
tk��x�M���P �:F�pq"���9cGL�m������pD�.�$����1Ȍc���/�%��d�PK� bʸ��C����3�A��"����7w�W�ǰ���J�b���u�y����.�*�=~ XK�O�����FX��H��4��n�e���ڴ�0���D�Jц ���/�b!'�۴e4z^gj�M�C��|�vP����T�jub��V�o��;��+"�$;���~�tW�	T��V����a��rQ�9"��I԰4��~��!�Xػ��A�h� �~
\ɠ>@�����l�>PE2��3g�h�EJd�|�����P@I�&/#��H���)�/bL����A#���O�����\ܔJ���ħQ�p���>A�\lP���ThL�ѯ�D��H]ڄ��d�|�t����ls?�O��V�7�O�������:Y���+� �b�1úQ��A���ۨߥ�CƆ���_���ǢgA��x�9�f#9(nt��au�� ��)�h� ��?�pvHh�
�ݓP��;L0�!����5��J1v��P����[�U/Z�f�N���~��,���PИy4z�/{����Y���������l�������Qڪ���4�N���vd�~Ga]nA����TK��-�ZB��1�;��1x6��z�k�u?�G�@+DǘKkm�O(�;��t��!��ʌ֏�6���ډ�Sc����Y_c˝�`d�h���������6�	����%
���^�G� ���F��
���=�HW�r���b9��%�q7H�>u&C��Y0�#���.3�&�im���w�|��h�x�<�6lqT+R޳���]��}P(�����#ST���標5�rh�WJ6� Md���
��:� �s4�lzsYWdVG�=4t����m����(*3m`�FF�g�yt*������ڄ�/��(
o~�a�b���3���~�ӹIoܶ�XO�'Γr���Kɐ=C�l�v�0b�g��U8]d��C.�Ii�L�(�գ��_+*�f�3I�]�y��Rhn��T���:�#"����!�²f=��O��h�=px�]�@h�nrQ�g�S>��Ǝv��꫋���7�@��`����tOy�U���^f�D��S��L�s�2 $�?��i�se@�gq�q��7�&� �U�i�$y�X��xR	�j�:l�>O66T�N��ORz�2�	�B*ׯr�T�܆E�B~K��<�z{j����ؠ掞����E#�'لbB���Ə��Ы��_Q��>�T�k��:`�A��亾�ﯟXΟR��?⬍��F���R��x����zy����MBD(����0��C�Ϙ& 6�b?�]�civ�5?c�IŴ�}p�`#}b,���i��N���A$KjQhH9�[0B��M۹���xձ|T�EY�{R�����`{y�br'u{��o��=���竽����ǫ�0�3�Oږ=���w�B&�Y��i_ōWH`J�����47��c2��hZ�"L��k�'���aB��!��n���	b��P�'~��fMְ"�����^�.��ր��i�j�Rup�Xc��OЪ��iT�6᭳]�d��@U~���	��/+G�D����/�oɜU+��&y�=�'�Y�$��V�1����wK�\�cXv�XNX2d�8��WY�l�o�#�ec�tr�N�gJ����}t�s�2�6�Jz,�
�1y7��S�2��W�!®�%l4����y4YyD�Um�ux�߳Z���Sc���!^��sV�?���E��h���g=j��,^�L��D����lI��qpY��(��$47�3�Y�S�U��2�.�x��E����9#�ɡ����%Lk�m$���:�=!��JԞ���F=���u��P5M���I�m�����I�1�=Y\W�]$�WxXle�?��6n�u���;=0J�<�ZkW�fܮ͆Ns��zT�:26�N���(}���/�B��|��J��}o��]��E'J��.k�}��s ���-�^Mwh<�7R�C��Е�[[�)a� ��l#Ї���h������8zIکXRT\̌�F����t[��r�p�(�g��'�g�p����6u��:y�����B�|�([��6�{9����#@q�K����p!4���N|%@��� ���ˈ�8�c�eX
�ऩ-ҺWa$�5�:���1�6�N%Gө�\f<��������n |�Z���45(YN�+���j��rG=��y��(ԭ��@-��P{��;z]0�A4����ۺ�t�v0��թ�p�Jdz{���TJ��-n�Bz�� �|�1"j����7�Skm�&+�ӎC��p��1 �-�Yҧ�@d5��1�o�,�/���$�I�e�li��J���"[���d�q��G<�n��{����{^rz���h<���;3Ѓ'�Ժ<�h��Z�[{��q�S����������7g�Ow����wY	��ȏ�'`���'�����0 �³oe��#>�d��R�"ɔg��F�p�
aTBͻǔ�,a���wh�����$�m_��`�ʥ�C��0��앤�����1!G޶����o�?j��J���Ѹ� o���$���Ǯ24�����|ԥ�j�3wS]`-wN�u����r$cЩ?�f&ʯY�p���Z1[Q��j�i���bT�vk��עmh�Tl�Q)���i��ѻ/:���i����s��i��a3�0���3�=.Ԗ��뉏1��G6Hcg�����s�tdz������CN�{�T�m�2�}����J�0�Mu�~<ص�B�mVu�W��~�Oj�Ȁ*]�۴#����\q��^g�j]�	�N٥Oh��ad��!e����d��+���M��\��$G{GB�.J�|�"�+�3�_R�Q���sKO�;�`�kJ"����u�O�c�ݶ2�{\[�ٴ�W�Gμ����}��w��S��y9<��j�.�K@��{m�������n�=����(<���CN=���U�eKi��h�Y���#3>��˳p���S��C�9�ꌪ�^��u�{��NM�'�J�_��m��(�d�J�:e�VLE�ϩ�ePܮ_��m���d��1]��)\���l�q��F-�F	l+���"�N�w01�F�����߫�l�;-��<P�r?.�0*�u;bVk��&��5oV5!��>]_�u��%����HSn<�`1U�E�?U����q�P�fg������A|���^����z��%jJ&,�Tz��uf�(��S��ʗE9ҕ��k	7�M+�`��}��uq��e�u�F��6�	�5���o���x�=E�swZSᱬ3$n�\����O
�t0�%ɔgj�7a��5SmBj(m���m�ƍ��p6��� }���?n1?���I��������I�(����}:���ѥ�U��)oJ���ق����#4I쭘���:ؗ��ࡅ/A,_T@z�Gq�e�o�x.���Q����=��nA�u���k]�AS�7�"�y7�¥ ��/I� ;n��o�p�M�,���F�@��OD+��
��f�@��w�JӅZ)~uQ�0g-�*��=W��Ġ[��B�x�o2ʚ�5�0]2�\�i�1�v���ݞ�)K��K&N�̄0�
g�����L�z(i���YG�
C�wS䝷;�!X���"=d�Ng�cay�����"ׂXf9e�cb�D7��KX=�����_b^��o�z#E䁭� �S���5Hj;�\Z¹ͺ	o8;��-x���������m]��:�ǁm��~s	F4$t��XOo��p�	:b|fI���7��B6o��2wR�২ʆb��W���ꬲ#c��YE��t���7��y�C�ջ"�F���%��T�F�ow0iN��/a�p��_�,v��^�/�h��4<�9/\1t��<�y7{ݭV)�b�3��_��/�wPv{���8t���y�@�nz�E �ҝ�,w�\�[˝�D�H���8�A��^y-D�T�r;�M= �K;��d�f͠(��n�ns���V������S|"K2l	�i3�f9��Q��ˆYT_8i��,��~�>^�D�G3��C���i��ioy(&���vAX"\�d�H��z�.n�9�E1�3���������o��k�@%��44��j�,��DTO��qF?���h���2Dh��+C�7Q��'W�nJ\�f�w�m���#�5�����r�-�#�ǹ3�_�Lȕ�-B�<�S'����K�S��bH�u�QS�� 	ܠ˽��m#��^�����̶�ç��j�=���(�M蹝(H�E�]�T��jz5t���#1^*ЊUMF�F��7�,�zdѺ�D'Aξt���^h/�y�Np�	�3�Ѻ;.�$w����[NHjһ۵���L��2J}�ˠy�/4I���S?�WE;��?E��oI'U�n�#ҁ��Z��"�B	����޹?8��t��{ў#T�ToҾ5*Q�΄Y��!`�'��V)&�a�F)�"/��l]W��uӺ�0�����3S*�bګ���] ���64�F�#%~�&> ����\��6+A>�k6�0�]vfQU��sP}�bupA�<}��8�O۝\���] �^�y�$�m���t�G\<������fp�"���T���d�P)0�M�#"���*٢nz:�J�� �D;�sy�� ��l\w�`H/rW�3ʬm���|חBK4�B/�@j��s�O�븰�����ti$���]~A�ޡ�`�1�����	6~ߖ��z�w>508k'�.�����h�@'酫�}��bDO<~�r����$�z��}���l�������W�Ԯýl�2�?M�%B=*��܌'���s��^|��E�4(C�Tc�{֞�c���o�F��94�K�&��Z�J���/�AĄ���D��0N*��k��{�JY�$^�7�j�*�'�`���	�7��X�#D���;�bG��)�ؽkISb���KC��yP�Sx*am����)�Дt)!�$*��rY��0�-dD�>31Z���|�����09ҬOWde]���8�����ly6%�#n3���H��F���b��J|	�o���>�����!1�賦���V�q��$��0�1�w�wl
��C����f��3�'�I=�#��X�h�=6y�>�l�S2|<��0�69d�}�k�$荻��D����f�1ąf�����4������w��BP��}���A��=n�� MZ�R�`7�J�)Q5�����Q�+$�8c�V�p���_�mm���ٮ�MZ��&m@v�z�L�N�,�k�o�K=��@��zꅭ�}�l�M���&����.w�v�2ġ�2B��{�E^y�Θ���{����l���:۪����{��>�����]���mbn%
Ld@�j�D���S�����k�x�ǐ���&��H�TL�/o�}	,���4ʬo���#L�F5�k'��kB��R���Z� >N�;8�����9��)�T^@
��ǀ��@�J��]-䫯�L˩H���I+u��2g�i������s�����-��)��
� [@���������VY,wgk
v�(N�O>>f��p;����V���=�<�7xO	91L��
o����J���V÷���NA��[�4(��@7E�`��sb�I� !��_��^��`Z�o%�w���(�ZQ�O���M�	�_�5V�w�|��+P��|��|о�ݛr�z��?����������Ͽ\����m�ܿ�z�|�6���!��`�]GMl�b�a�^Z���^�KM	���f��^#4}�;^yD0e4]��ւ��D�љBr�`�2��5~�)����ufK܃v0�Q2���A��Qg�F������oC!���ݴ{��}��VI@��-��{r��\X��3�0E^f)0j�{��un0!�����V^�o�\a��6c�?/8���Z��9WT��˯�uI��0��5���*8fHbg���@���^�c9G�#>�a�@HA>F,�2t�8[#E�H�����Ϟa�pV}*���C�:��r3�U�e�Rr�ߦ`�U���� ���QJ�
�<'Ǘ�i�V�ﮭa�nK�Rn;�2�{Zbݗ)�7�dl��!��N9$j�L�?*?���d��m0�A+�o��uY�t���&ԕQ��~P<��-J�	d�5[��<���EU������X��JT�����47�JK�QY&NRI�ĵ4�8�-��X�y���������g��)�M
:~y��|@� ��y����߻�C.N�ď��4����A+�������q�Y�Ё�tZ�״���Ai��w`A)zp�%� �#͡��x��Z�	���$~N���o5�̂�y�[��7,#������6�?�n�Ď�h3�AW%f�,��z�쐥���[�2F+R0��E�w#c��&��pc*�Y�D���﫽�_�Jɥ=�~���ڕ���;�S��ao�GHE	Z��x~�o<(G�8==�F2Z��7X�i�;@��mV�$�t��n1���(��H�y�qc�MH�X���A����(���C+=��f��,g�s�@x�2]��{>��zG'�6h5���LS�."z�$�n�l؞��Zط2��n�Y���ܡD#
��������	��]��\g��`H
�-��U[��V������X�����bR� _+%$:k3�&��9 �L<[�G6I�XWq��,t~�.AU�%/D@XF'���MT�����8�`^F$M��l5.�sA��:Ph3�����44����b/g�C+ �}�<�]��Q*���fu�E��A<K��C�Rc'��⣆P�c�,�
� ���tQ�����S�O��,�c�C�e�z�0(������J�̃�>3�}��$�]`ڌI�� � �8/j|���6V7�g*���Q˽�n�g�9���~�;^9D�ݠ#VO����fGKN�u�jԪ�.����ꢚЕ_P���x��x��~�֫�-�6I/�b�s��yH���1��5}���5��1c�/
#v��oh�1p��{�Ҙ��4��	>c��<���k��u&�@�����V��\��=�bm�D��4�¡�`�����Q������
�c�o����{�˱��v�}�Q5��R�x�i_&M5�R��Ԗn?�sL������|��9����Mo��_����	fXSoM	��thi��p�~�4V����܂����7�_Hi�#|P�ŉh���J�ﶪ��_3������T�f@Mw%@��e5�&����g�CL`�y��@��WK�&�9���;�����|����  �4��c���_]g���r�CS�X�>���F/��k�p�#��z>}��K_��1��Y�!H7�Y�K��_�TW��nQ��d���47�sI��4{H�H_� ������oAz^���B&]˂ ���)��ʗ)����;e֗	Z�𣁞Qý7Ӣ-ob�q88� ���*
�/�`���T��A`w*j�u���Nm1��6�[�t7�Y<��oÓ�>�/�L�=����Y��� !�e*�[�Y�=�K�d���h*7��&�����a�1&Fq���61b��ٔ N2�4@Mk�fS���oT����;޴a��+�m\c2*��qj3�A6���李z�[�2�����D:��[����)a~Ё��e J	�E@�}�JC�����-c���"
�qx'>[4&���?A�}*�v�w�>"j�㙁F�EaH���5�$���pUg|�Pdc#�?��&���0�!�v�V��̄~�[�_a�&ci57*ٗ۲ڷ'�;��Wéߑ�	�T������I�Z6'M���#�;#Bv��l�닌�s͉`h<�B�� �9�є��F��لV�%Y��h��~3���#w�ZxwvÝ4�҉�ȹ��5�Y�>��P�!����]�9�,f�Jwz˘3�췧l�ʜ�L#9<��=��v>���>R��y�0b�߯ lJ�1�Ҷ���*M:���c�B�'� �޳��*� �h̬��S�Y�j|y~��_?��Y��6�Yb#w[��Cl������E��ꪑc�:��L�ʽ�AL�����,9r�2�����"N���hs'Gd��͗F����� 	Ր���b-�����\�h^����^Zw������,|��դ��5ַ�y�?��NYDo�v4G���� ��&��}���e���'X�Ptgk��?7�3-��m�k�.C�O�dFޔ�PfƉ�q\����PȢRpfs+s^u
��N�;�V�t<�C�/��b�2�'��\��r�9C�Y�C]��L1H.�	]�9���ʗ�jV8#aX��E7B�ty��70M����{������?����iA�Vʂ���	HR��R�3���R�����y<	���@��_7��;_��h�EG��������U��5b�,L���[�*?�z��Di��Y���ݑ� kF�l^�81���˘�3��\��&����t��^L-��yc���8$���4��L�	ۊ� $�("������d�k�!��B?Q����lE	3�����,,n$
M�qF�����U᪛ߍE�n�t���G���JW�`ņ�q�*"�g{L�wRʩN�}F�����H5@dN�A�wB��gk���;И�bB%A��nb�7����;}�tFQ+!�U�E���wT��Fo�Ք���0iDő������n�j�
Z��$�������|w/�=�<m(���A9j�b�9}.��-ΰ�ٓ�>&��)��Kܻ|�������b�(�$V`	J<R����fX�ux�Ź���j��s����x3��_�a��,t�u�j�3�6.���2��uҝ�tikZ�m�?��u�EN�hhHnU�3�r��3
��z�	�=�2���x��z�d	�ϮŇ��W*���Q��vq
<�me�v�t�Q��ݗV����]e��@	|l�S|�@z^�Y
����`
���6Cl>�3RH�{mph����mvwA�� ����"���s��0O�Y'�m'ܤ2_ņ�O)0�j�Q\�l<A	�7e<+����/��t�������j�+ׅlє��򲵸	�qފ 迚f��¾�I�r�]=���"�T�<0�ĵyͶR���X��@��_E�+I�s����xFh�e�{��F����&8�Y�����6�ϴj��U^?`9��֌�Y�ӑ�x������]s�w	�y6hj5I�p�����Ƿ(���h=&����G���N�����tUT��ݼ?L���GuL Ns���J~>0�f��;5MAm�ɫ4�]6Tl�p
R���2�4/õ'ڢJ��uc�ę�sy_��ɕ~�`��������k'tR?s��a ��V���$��D���� �����W��
��Z���bY�>KA�^J��n�LF��PC&&:3��S��~�E^�%��E0�f�� k1�@��c��'�q{����@��}..k�^����vI��NuF㫍��(
�Ӄ�6]j�%RN;��#��s�P`ti���f�~T��L�%�9�9p�	'��؃���Ga���٥���kI;�&�����Q`��y��f�&bC�3N�w�8#ƺD�?lZ���c�w�$��8�����
r㬷+�'������Vv͔86*J2�XX~����d3ʊ۰�}��:3|��D��Ռg3�c}��QY�6�|�3������l��2rG��g�ܦZ���E�=��Fw��[��)� �˂�KhCM�u�e��x���ؤ�OM�� y�_+�@O0庺n�q��%��"�Cf��M��s[Wkm1oFn���Ц**���?+
q�,�ub#���2�l�����vt��;��6�DLD��g{(��_�*��_^�e ��-�p�s�����G8%^>��]��������p��-��YǳD���F>W�ew�@�}�9�|�O�	Tq�Mōs$���2�h$���^Pw��
�r���M��^Y�y���3�.�w���ۚ;�>>���k��R�Fd@�VĽ��.x��b䠀M	c��:�� *!�4��{v�TW�(��v������o_}�Po��͊l0<�gٓ˶�Ik\���$(/�2ԠC$^!~&e��A
xtE����?@iL��;��H�y����h����Vt�}ɲ�4#F�7Y<Z���P�`�j�(��M�Z��:�}����hΥ�t�48�/�� �����UYdY���� �Y�޼�&�p�gV��� �4�B+-��asU�#�aJ���7����ɜ�����h8Y�IdPr���Y��LF�♠�HL��wP��<��}��Ѯ���*���#c��.�F���;���v����ɟa�=¦t�D�_�qx�/�0X�pi��z�w���|��o6o�þ�l��D��i��%�g[д<�� r[�IT<H��r#w@G!V�o�o�Im�#���ن�A�*�^nHjB�
8�PO����r2A�b�odSxJW��[�2����g��m�_�Yd^�"z��=�I�Ar���d�_9Xu1��
	��ù��0���v��7^��.�p�������.N=ew���UѼ �ۻ�����5N�ސԞF�W8I�s�7������dxÃ!�7ŷa�Jt��t��H��4AW�1(�=Q�;mvfo�g<1�K���	���r-V��ْ�`AN�D���mQ^7u�z����3׼�v5=�C����0�|��׺X!�L�����P�9Na��0z%��p_h~W�N�_<c�	1�pAt�^�Y']�F�P�=00M���2���6�E�����,�x��=N�o}3*�<]���oIN���4�T;w^�{�g���+�KE��׀d@�������IXWl�L[��qu�z��
E��]r.CIa���l7d2�/D���@7��˹|�}#�O��B�*°luv����;�@4�J�$&͙��D$*s�%&���fK..�ڲ��x����ͯ����L-~	�Z0 jh�������'��=�ƕ8��,���)�0;=5[�k6+�9\
�]�ij��Љ���%�ˍ�FW�Ή�6��>�B�^�`��F��������3�V&7>w�}$��ES���ݩ�Ɯ,R�U�0�h�C�@e#��/�-��h����0������TV���7F�VV�`%;5g���@i�"�8�5ށ�+T� �tnn�6^���t�rʆs�F��\�BC�n�(::�/����L@�a���O�|_ɰ�['�S�!҈��[`��ʴO7~SVD�E:�u��u�)�U�q�����	�v�`#Ts�������>��TU5��qxж�e@���#��1��js��Y<�6��5T�y�.UƂ��[�aeJCt�^`��׼�S����=7�6�z�Gĩ8�f�s��wnM����x����*�s[mv��J�d��"�Q��x��h1ڌ&��kWo�jj2��/Ga
$?�6h��ݏ2��*�#$w��.E-n�L��H@�
��vz�T�g�FmQ�dxT}#S#�'��mY�{~x�� �i��J���^f_�s�B����&��v�s0G����03�_�?��4s��� 
���V$���A6? z�ČdX�5��*�o���[d�'_6��n�����2C�1G���O&.�w��	��`RX!�"~f�;o�F�b��_t坲�+�:/6%i�~@�n�{�EFǈc���w�w%�TJ�xn`�H1r��|/Kk����l�uL����T/7�/��l\Wd�KQЮ]���I����,�*/R}i�?~����.�%�"�l�u�;���:���%Z���`���b��u���3ϳ ;�����Ǹ���-�P�H�!�{���l\"�\z/R�ǥ)@R��s���f���W
��>���x�M��<�*�f3^��������h��ԑy�_$׾S '���DT�S��� #Wl�G�Ukͧm��r��s'�P	�h�)�0I��R�3�7��P�)�]m���ڕ��,�$���?dS���:�P�����Q�����X�"F�蟫|�?��"�)�.o5�j5w���k�4��ϔ� �i�֡��P���,�yV�t�,�i�^dB��@S�O/'�"(���@���o����VkY������s�G��D���Q��,�Ӷ�I�}��=�˄���:W%D���n�_�L�6�fX_���ڽ?_n�S�By#�3�JK�DQ04i�v�UZ��i�eH*a�^L�ya*#����P��7�s���XJ���:I ?��g�A��	��U�M L�5�K��3@��A����b�e�}'`���w�S��菺�R^Mj��әu) �\�T�b�b�'���c��q�����Ҽ�ժz��X(���L��af=�(l�>�����x�͝��Fr��r����Ju�Lܢj�N��b�= ��=(�طv\v�Fw[�:9���S�jQԒz*0�XEC��୔.�7�o?Xã��+�
�k1��>P2���{$#q�QQ��2���g��������;�214�9R�b!Cs�'�H�'�a���ݸy(��0�	>fb�r������~���+���'k��wF�9��/ޖ��V{�͋p�d��I��*������@b ��Ø���I���Yr�ߪ���BM
�G'���+q�o�=P�H!�"�����<z ���j�:�	��d݃9��;���?2α�>֒��4X�ԛ�^⯈���:��ݶG���P\����U1+.j��|A�H@A�d/��C�ar��<h�	 �x����B���@\3�����������$��2���IL�I���Z".���P��,"�zN"�|{�~D���@��@eDp� |p��g���,?�� ��j�T�ه�(M��Ǔ�jk�O|;k���9�7�𩈭#8=ฮ*�2a'����強&d�x�z(	�>|D���m��]e�H�$(d�7�
�e��^�fj�Hn�� :�x#y�n?7�Rs²�a�v�6bY�_��`��W�s/c��{8�v�m �;����U�~�|r�h���o�ñ��������;%� 3yF~n͐���*KuO"m�ouPSw`e��d��1�>d�t�WT����oBo�F��zNvV�,e �~����8�3�n�����W���Zd�Ob���\ǮG�JOk���3��`�AƎ�+��W�CVtU��]M�v��>,6�3�=�[�怭0�V\V"d��4�re��4)pf��lV$��z���C��$�)�Nx�{��eڧ���R�n,6���:�L ��)��N��B	�����壁����*�{-�C?��$d�����f����S�~HkRhtR�\'�ʬ��Я�������������9JI�]�Í"!�˺�ua���� ݝt�Kj�H�R\�!%���X��s���'��ģQߙKf��jC�֎��@=cH�)�3
I������["o	���ge�0%��p�#H�"��;L&��c��Q���m�E��R��U�H^CB���p���w#�ź<��?;�|�fҠ�w�!f�t?�o�V4��$~��.�JC���8��A��ň1�{�KZ�0���N���4�:b��D����#\ҹ�k���L>kQ���S��B����9
��-P�ҁ�9u�����6l+�c=!U�̸+�+L���S=��׽Ʉ��l����ج0`�`(��gf�<�D���k)ݬ~GsA���䙥/P�J�'.e�A.I�ǥ��!���F:�1Y\��!�
�$��,5
����;��Fo�/�|����O~�ˆN=D��OWH����nt]���A�fGR~���g���^��_�ɪ�*��C�F�#��q����&0�Vui�z�o��YO}����Y�����x?	e�-p1���U�E���F��@�=�V�
\3e��ⲣ:�;��Z��a1��~�W�ojn j�N�Oᅔ	��Ðl���y�Pł�D��>Q���1��/.�M�-Z���+��x�x����z��s�!-���l��DI��|/����ݭ��>��i$�����%� �D3'��* ��4����᰿���f����Z��W�������o�lK{Gd�U��	����ZqV�h曧��}K�a�-}�3��; e�4���f��3���UuV�e��uS�EL/@[���[��1����A8	$���~2]�֯w����=`�䦆Av�K>yљc�L�e(g�9�b���Pk��9_��QB�a:҆&'5IR���]Y�;���	Z��_�Ky����VI `��L+�8H+���ކw�?!)��~�L(��;���YiEnX�{%��@��j���)����B����\HnO�4.
��A�������:[L��0��.4�;y�>Z��[���x�]���3	=K#�/4�?l�qhM̱���<ц�`����#�����=��^R� Ўэ�)�@���2�=�H�.��[P��)#�%i1�U,֖��T$�mXk��]���Z���XQrd��
/���R�!�<���ndO�	7q��]nd�
��7NrCW?i\߲�(�슚��r;����8s+[�9	��SC˝�q93}it*ťž��B���7KN�ğ���G�Y�3�}g+��F~���U|틌���h�m���)�?�?z4���e�����D@t�x�7C����&ܕ�hp8��q,a	"�",�Q�N�� B�`@������`��ף�T��m+i�0�)��jba��4�1�|.KX���ng���C��W��J��m��F�k��8(;�L�|ϽsC��4�w�}w�&��,Rɧ�ߤ�X"���X=Ĥ���<��*�=���P]h�ҋ�=@�c=X����������=+��j��1!5�z�o��:�^T�t7		���;RM[M�<a7Ɍ�&�锺T��[%�m.e���U��&6���΅&���ϯ�f����إ��/h�rO��>�����ND����/�+�����M�qrS3���'�p9Ԗ��<�;%�{#
���(�-�^��S�J��sǥʷ���۷ǳ:��죫�'Q��zG�%i���{��m�р�V�x�6�+ԥ&���j]A��v���L�}4�!,b,��ün�ؔ���)G��N��X�Bk��"[�ݯ�l�!���Knu(�-�$%tٽ^!���\�L�?eύk��O	%��-�'s�@��Ζ����ʹ]�7������оv�(�Z+����kѣ�U��bOs�6q��� #}d+�Dl;M�3|Q����+�dI��f�_m��"�m����1��\LWt�2��#�L��*te�(��n'"�f�V%B�M�ޠ�Qc�bcǎ:m��#�˹���EB���������oi���w���n�L������������X�c�N��it���\F7��>��ø�t��˗�Z�=�V8ʩ�X1Z����uT����f�YNp�ԳH͠��(�;��XmGdQK�Ie�kC��dl>��d�L�q�'���H�PAc�	;�@������uѪ�.Bl(+�S�=��	 gCQ��ƲT\��� Q��L
��<G�mi�|w:'O�ތ��~2�j��F���"-�Z��K�9���e�ǒE�"T�M �D���>!a$ .�=%%h ��e�
W]#�|QU��H�q���3�₍Ge�v���ך-<s�G��(1���K���3O�E]n�4P?��]���A\@g��� ЀY�$y�Џ�vH�(W_��}@�x��%�ޝu^oH� �om4�b��w��\C���%�ӄY��X~�y��RX�$FhV�i�������%��h����t��xԫD��V���LZn+P�\�0%z]#�ũ�|I�8y��j�
�KsE�
�==��}w�;V�����Q���a�N(0������c�n����g�0_�;Q�@��p���T�o(ɮ�F��[�)M	x_���4�R���v����$OH����F9WR]�5���p��j�M�C;�fdbC���?���Kkm�y��1a���)詤�&6�$�?��R��-����6���<��hPF;}c��v_WQNT�@Rw�T`>�L:����7 ��E���쀁1Nq��^u��k�� 34��۳(S����Ԩ ��E�@���/������i�'�)��d��"�G� �|�&���<�R���;�7y�
��J��o�y3۶�Эˏ�#����IŸ3an�@�+�;�5�i�3��Ǘ�2���˱=9�[��_H��Sqv�௼L	hEK譂�/"�,�\� �@ =��7�)�{'I��4�(Aɶ���]D{:�KfM��� �y�i�'���e6OCit�}
��tv5�$�zʿQSz�(J΅\x�;݉��%1R2g�ke���>P�zQ��XErѳ��+������D�������p=��g0EZ�6�>o���)�h+nci�Lz�B�\�#�ᇇ�HfcS|��������n �X�Ъ���VzgI����`�ԣM�p���w��h����|�����:��߷��·uCo"�P���:�#BjDЅΜ嗂��͉���:u^#[�Q"�{GG��s��
��U��Z�"��ݽZХ&��Y4na��p=��K�$Β�����ZR�j�׬��[=�$�0�B+��L#;i
tޥ��r��3�:x��la�y���}�����)>tJ�j����NG|��'~���%��KMA���G�O��d����㌽�<��*'0.�cu3��D;~����\���O�e���� [��K/>T�R'�H�Y�o:s��־¢5����1x�`e�P�g��v2]8=\�q�A�������|FKrs*�ʊæ�2�P�f�H�lڵ��<��l}���2}>�ڦ�b����F4g�DO�E_��`�E��w�ҁ��c�e���� p�+T��M=����TX�R��W:*�7�S�� \����Eg0��i>��a�ඏ�Uߎ05ؽ���ֲn��E?А�v�g�o
љ������ą�肅�F�[%�z�PK��1MIb�*�GQ��0���%�H˼�l��Π�͔� �|h�ؑ�,%�?Ɉ����|iͶu���q�6���ܶ���\ܨ$h������c��8���+��e�,]}`Б��x������'�E�����8�Ut��CG>�<JD~���~�P"瑼Ե�,�DZg�>�C$>^;�����G�B���di,��uۮ�!�������7/Ao��`�!>�Ū���H��E����m:��GgZ��"�7�n��b��
4.����t�0��IR�����ޘŨ����q~�F�K�H�T^����+���ۜ�6B���8k�K�>��޼׵~�$6�T�_ʶ�"�P#�s��3����Gx>@�C�!��v��l8�ZۉFO&#u��/�Q%�ʾ<����X�I$���,�38ؼ�NKΔx(Q�?�M x��:�r�pI2��Wn�C��/L�L������Vm�8�B&���ڴ�m1@=r�,��L{��������iܠ�^J$��+qt,1O)�crc]�]�rբŊv)UZ4���t����cC��x1`f͏�k�U�����$蓢�����6Yg&�H�U/,Nа�4<˸߯m�#e�4��6�3�B��'Gl�3ۏP9%ٸ�X��r�:�����+(Τ��(�|�7���R5����;`�b<G�� �a���#��p|*�>��C��7��XM��$��˃ޛ����~-Q8����
#�%=
�0T4,&�5�;^@��Y�6��Q$�3^T,�.�i&�ҭ��$�(�[�y�[��{i�^���������X�T����8����h:F�q�e����+�b�y�*Kw��6�t%VԀ��izЭY�@/)m2��,�Y�q�������i4�n3�I�h`ҡ�7-�t�� p�1HF�^l�)2�!�CL���TND�t����������`6f~$��t���f>C����4�D�ɯ�a�g�������o9Re�`0#�so�{�h>.��m	\�*�ţ�Ĉ.%o�����0�?�$������K��J���Q����/%�#
��ՙ����m���)򸡼���*>j�m\g-�d~1]4�����jS��G3A�Mυ��U1�%��I���|���kԷ[��l�UY�E�HÞi�R����ؒ�M�>!���6���M�o���^
����&�="�#�J���;�D�U������4d�	���u�G�[���6G��D!C�exQV���8ҥx &��
�]��=��ܝ��^^����ȇ@TDalmn��K�ѳ���<�j�(��}�v DW_5�3FV! �9 Aڣ����6�
c2�-�o������u�2xB����{+E�,�b_Ե�	��9�-?��_+*mTTj��i>s�z ��
��*��K��93���^E��u#�@�M\��m"a��|l�~��
E�*b�:�ׯ0E�f�[�JD���f.�m>auF�G��c�ņ�q��<N��V�B\�Fy)n��!X)��%�
(����JZ�"ރ7{�1��6/���c�&���/��72e[C�ݸx3�$w%}d�*ث7o�>#��>�fK�L_ڗ��mL���@�t�������WqR�!��Ԝ��YP%V�p5���,}K *]��Y��� 1��_#��`Ҿ�y E$��ѥ~���s=:�b��O-�.Ӣ�+�����&�'�L��x��!_�*Q���q)���*F��F��b&��<H4�����a�=�����*L�j��*R��F�,�,�b�<��ak�E�� ��v�2;}�����:5��n�KE
Z�Q��]�b�Vn�@TD�E������q�y��H�&�;+AHv>R۱7Rt"����pab�!�,	�w��u���r�wA�,�uoѐ�D#�0ǆv�^�%W#���y��S]L\vŒ��B��/wŝq��wX1k����bf� �����!�sӎ��G! ���KI5Vw��8��� �A<���`����D����nK�4��`jI)O�"�;�}���J��aL�{�T<���ccR�B��Yn ̃�{h�2�mt��g��2x;~��%k0v��V�<�d��]|,n�ܗ���7���b����:�Q�50�xX�c`���3������݋�r��|}5+&��N���臒0u��cR��&ѹb{J�W���`P��CH
�=O}���m�~I�ҫl�W|Tl���_0��2�l�`�_?��Y��2�Q~�}�Lb�@�9=:�|ʼ�W.�`����D˔]`��L����hu��o���|%sb�Á�h��lA���bIj|A\�x��������2Sˁ7g\��]��|!VY�%o�M�c�
�N���C���G�+=���$aA���WS1.�}�'�+U�*��FP�Ct�M��z(+I�7f<;<��B�//��^�+�K/eo�u%]��亍��d���͚5~s@���|�!%]a�l����_LWG�Ȳ��0�2S�[�B�dt�`ttѫ�P�q�DQ<Aۅ-h�2��m����{��K|���ki�S�8�x��׽��+M	��	Em ��X�6 ND�}�Y����k�|&�
�[�n/��n��w��X��Ӈ'�s��/�@H$=��Q�x�q�o:�eT'�l������2�gc��42�-g���n.��9#�O����z���PQ7�w�����J�Pa���'Y����m�0���bT�Zܫ_��@=������$��g.b��<b�vscb5p��:�+O@��ߞA}���d�YYC����K����l���=�x��kP*i�J\��ON�x\P�C��C9�נz������OX`���\F��V��2��x����b��&-;��W��%�3
K�="���4i���:k�.Je��'_Xt�Y�p���vi��V�4mW�_,t >�^}-
<�Wv��6bG,�\n��	��tB��囄�[�f������	���a�� 2��q,�'���턭:��}	�� ���Ssh	_ڿQ��/FH b%TT�Y�A^-�G�躆������:��J�9��%�sdK��	�I1X]f�i<V�
��(gu	�
����[�E���F�&�΅Zһov�J�87&*���H
[d�16_�!���r^t�X�{z,6yx+r�6�-�fN�lxf+/�hOP�IeY����f`<FṕJ�z�g�5���fv��-����Z-����K
������C�kTjq�p���D��X&5���Μ�ǚ��"t�<���b�*��Kx�� (e�1�ޏx!SN�7Խ"S��tԼ@�Z§�lؽ��� 8���P�c�󼂟㖀5eNc����B+ƶZ�( E �ztN���/0`�f�B�:JP8��2^ɾd�>Ϭ��qfIxm�M�ۗ+��f��N�;/跘�y&6RS�8�&�&I��i�\�(p)���3N{G�c'�1�HH��C�I�v��':p7 �9vm�U���|�K�.�O���g����qn���;�c
��LԢ�,4f���9�5�l��f�F����U��^�������U{��D��,:Ö��i�ژG�ʽO:�b&��)���}�c����~���z��x �d^U�@-��[�ث�~�X���<�7G��&b�1S�� Q )��� T�����-J��I\�.u�e�� �C�앾��w�`F�g�0��o���lC�˶��*qr���U�*R�e9m*j��p�l*i��!�f�e�[�`��!�'����E�n�)�d�˵�&�J��j���`;Y�#�C!�_չ��_8?X$�*@�Odю��\;�@���
6j�6��NN�!�­s�*ܶ]�g�?�j�ř,wڼ�@���3�O,���+���"��C��5Z�}�6�/z��G���sHjn�[�Kɚ��%!#@6a�s���C���譑'�}����GԶǤʒ����/�c5%�EM�L'&l���3�k�g�֚�<�Uד#����j���Rj܃��뭔��p��1�k8�s�������bm��S���͎)�j�uɨte�G��ۯD��$��j�]��s_�w'��m�'�D8���ݡ�� Y>JW����hb��s�7�7#�
N��LqM� d�U�A�},�x}�zf^�����n�X�ݯ ��`vr�PB�0?K���|�ץ�Zy���*��5U�O�4h��se�V�,��D�1�>Ig���>}���z�y\�qM����o�-JhV6�8�I�N�,=Ԉc8e��t�SW�B^���:u�NAӜ��K-�z��q���K��/�nۃ�?<^�a����u.��9� +J8���?����%g�z���֧:fX̎=�g��F����ؔ��%}�.:dD����bɬA��|�ռcx�}���H�nEO���#n�8��������J�;�,2Py�;q-M�F�ꈊD�����Y3���1�����w�_z��8H~��@�|Y��P
��j�������P�Y���\���^IA�;"&�ol��l����G�;?���{mJrsd�_!�W����c�皝����"�����s9v�Z��o�3w����!U���Z�鐍N��T���>}eh�q�D}D�kv�}s�T�����͆D�3�z�켐q�,���v!}3��'�֪��r�b�uҳW� ���܎H젍��h���+�ޏ�,�o9r�}��Z6߾;G�ڽh��L���X�D~�g$�L�MC�������^�͡���焙�9e#�Fq]�L���&�PA��KF"&y����� o9�Jk��-�((���B^g�%�D>wY��ib&� gj�]��F�?G�P����X�|��k��9������V�9$������3e1�Ah{�m�i���z̒-|�ڷE�u�e���.�:�lN�R���U�V�G<�e�pB����!b���|�:����ѬܛN?\<��qp��%���k����^4E��,�vi
r^�,E�j��&V�/T.nG�D v�Vi�6i����	6m���8�n.e ��w}TS�)��
�Un��p1��9͏>�O��sv�i�ál�
���ƿ�	�8��2���;���9��"�(�ٗ�
 ��T�΁��S/.�e;$7�(B��2.C%�+8���ST��M֨^q��X��M���>ʬ�%M�@5?�3o������>6���6�I�<��=��67�j2�ZѮ�P����qG�fb���t��q`�\i��
gB����s�J��2-a��b%,2��\��SԈi~2JJ���L4G	��:@'� ��r�}C�˽0.�l\�!�ZB;ڄ�C�o��u���A��������$�8E�7�-���PN���My������x�V���׻ q��N��B���_��ƈ��k�>�K"Z��<"{�*����������ݨ���}�\bx��_�L�I��g��=�?�=�Y^	&Y����������x���!�:;��Y��!'����c!j*��bTZ����L]�2v���,�W���C�K��r%)�C�-��a��H	h�dk���yG���e�@�/�4��fYq��s�9�<��EӳV����� ɭׇo}��/>����gy���� ��t��q�V���1k��4�D4Μ*�u�w�X����0��Ţ
�}8���=;��Q&�$�h��ɂ��gA1���wF�M�I��,~-׆]�m1!���ñ*��Ӌ��L{�8D��ζc'������P1�-�K�/�^Iq��UΖ�ٽ���E3�h���3Aھ��u�!��� 0�?��z��Ĳ�u�/�8᳍��� �H,�;�n'��1l��_�ѽp8��>�I�q36��,MZb��&i#��Z�ֱ�, ���(���z����'o�B+'Ch��h�܄�2O�-c�P����{�B�n��Z�wIY��o��q����U���p��̼� ��;�]��މ?���y�޻��=.L �!��5
��dz{�8��ɝ�A稔�"�������Թ�sP�Y!C��:����Ipڲp�Y_�r:i�U �"���y�v�!!�B�t�J��z2F�NXbz��4��iR28�(ĦJ�!P����K���J�78+��u{AK���ς����eX��L2��C^��/9l���}���TE��ab`ƖuX�	��Q�D��J���c��{c�뜲��Z�n���Y�#� :2x�W�ab����	�B�ͱ��p�O47�ֆ�JD��y{v� ��9��{�B�\��RE�F�;*�h�&U��M#k��'[��72]�ΎA*�m<�7� Q��Y�yz�p���0T$�6Y(���+!	�rP����:tGI��c,}Ӓ��AJu��������Ѩ�b�6Q�<`�h�QL�p���O!�D�<�7��\)a��;�yX���b885?6� ���c.�.k4T�ݾ�)V�s���	�n�{MT���bq��x*�o��A͆	�~?5��v��^�T�����N�o�1q��?�+�g��~xt����G
F��K��+�涘�Jk9�� �W�K��/��jn�w�\�,$ª��R�jj&��ʫI�( A-�>�|z��2�H2�4�*`E����{y���<M0�a�	p@x�\�՚��p��ZH+Pze��^�A)���ӳ��SRW���3�U�g�ŉ4��,Xw3,�52ɓ�蒮�5n�����-�7�4��{S�w��9�
 �\��$�5u�ǟgd౺T��
��ݼR����Viǳ��j���f)��S��d�㜢��F=�}ٹ�
��ԇ�w훠�)�*Ƞ������p_�]/�T���#������|�sC�6n�L�9X8z%]�^���S!���5}hV"�UJ;�n����o#q��� ���o(�5��4|	������1y��23�<?�G鄂�]�a��>�^�[� �*O�"C~�Nl�U� �Ah}ܙ����w�j���	E�� �j�İd��wƆ'����T��D"�!{�tOýO�����TX�T��;�k��0�Jz#���g��v�Ki����6����7�����0姓k{T[1���bY��&K���$'/��E��]z�dli?�dM�Co�4�C���Q�Ǜ��k�\p�J�1犝H�}MrRm�M�lMqMްI��2 ��e���`�qh�P�A�Ga �rNn��S�F�������R�w��$0�/�4�;x�	\hѝ����)L����%:̟��*G��4�2&Z�<�2:tŶ���M6X��^Ch@g=<�t�|e����3dƲ
�����F�߂{T�w�h O"�-{�`�4md�Vt��~`�9 0�n����>�^��5�S��-d��ӧ	1�ަ�L�Ĺ/Xq]Kऽc����Y�?��Q��|m�[�� ��އ��E�4�)�b�^L��A��R�l������c�Ѹ�R�pYM0�Է1*'��f0�����*W�?Fy����[gZN��ƿg�jh�p�{Xl�C�P�M�r>�k4�d���W|���d_7SFj-h-���X�Mw���}�!�$���_b�k<e�AdX�ۧ];{t��m6e�`���7%��"�j�M��@xf*r�v�c2�TSE�~N�#!���Y�NWJ!	�8��p��y��8�s���쑀@u_��\�j��8��0�����W�<�������K���x�����ެ��rUmkT��acgg�@�P���_���Lz ��T����d��i����ܺ�{r�*]�Z��Xp"5j	�¿S�v�x�8A���<V�� �#+$c�V-�Z�oj��,� � =�;�!tbxO�G��Ru�R7��E�Jm�����_U�D�!�a�L�o���iV��I=q3Z�w�ج�-u7�![ԛ�	ܧQ����P��K��X�������`:��c�&{6?tq��IY�k��a6A��gg�	��bNo�� ����پ�8�8�>�d�Hi\�����LG&���p�uJ�a
E�bU5p�Z:�3�3����J��I�kE!h"�f�5	!w�q��K�8��˔���]��COJ7YEBu�cP�RԒ���A�m1�͂Czh�n��΁ݓ���;���e����w6*09�]���9��E�L�T�}w8+���7s�WP2дQ�K�2�oj�C��*ܟ��Cǖ���yr�u��@���t�Z5��=.�V�(�(���	����Ĉ�)���[�
��6hӟ���i�p֝㌁g������8��'�O�5g�C"�����@!��F/u���.~\�42xŁ������ص.zy+��cW��A0�r1"�`��c׬�=l>��׃�\s v���z��ѕ�&��J���`��z�w_}�5�L��j�_�
M-�6N�=Ij��}����Pq ���-�k8 m�;��ls��j�.���ߓ�Ç٬{M3^x5�0%����jB��J���Yޟ�"I��g���f�^�+��-�]cC.���	������hV>�`|H+���`��� ɞ��)|D Y����y�y��豸g`���8��J�7,�G�O��&Ɗ�ֿ���!=<b+�q?ml_���)�QV�a����x�}wT[]&� ��|Q_f@z���1�w��� �5tX���RM��aY����y�f,4?B�O'�V��TL�h������ѰӨ˟�K��^�c�<�ʎj�iD��7;��?�Hϴ�ڪ���2�bu�SA}���	1T�1e��_ളc߳�!j���ޛ�� ~�	٤L����,t��B����d�wWL,����]4 �R��_ڪ8��_�`��Xn��"ԯ��`1���B|Ӆ~ئ@�ַxT��b͑���r]��+�H��b�aQu�kJ�+��;H��������|P��������t4'T�a�=�w�(�+�U�J�eO�����0Pm���V�D���x���m���9�Ӕ���d�+�w6�\��J��rVs���>?� S�j�1�0q.R��H]McnB���U��)q�xh�h����{'�S�B��zo�R*9��y(|c���Os(Rs!FH"��*+��NJ�� ���@%���� "��#ˎ6'�!�3͗D{�澋F?���ߠ����i�>g���^�y�����G�x����}1ꨉ��b�]h*�yw�y~B\8 ��^D7e�Kξ��4��\B) 8�&Pb	�>d��;h;*�zO䶡qF,*��}���ou j�*�h�(�X�?㐮�y�_�_ܡ��PL�h<H������'�y��JE�`����˔��]�V��Y��$L%��n�s�3桾�h��Ki�6ʏ)�����4��}�!�Gv���r5H0���a
�N_����l?��Hc�k��dPfS쩽���KY��]�@i̼��l�dW0����\P�<���o��G����.�2��}���S�:]��w2�����Le.[� �--?B$��o�!9���)'�K�1�Tܲ��]���oX���J�,IcK��ʀ>GJL�!�3�,E]�Ծ]�~�&(��>����J_��L?/�⌭�%5�Ǔ+�6b�I�)Ɠ%��B\�@�����mw��x拻!��Mwn�RZ"����AhlHr2�U��N^�<�e���)�V��4v}�����U��%�i�����2���$n&�nF��'I[�GN��=�%�K]�keM�ٗF�,2f�h2&A��[�1Wd��j$t��'�1؎4�Ϫ�FTԺ������h��� �ܚ��J5dA��i��Q[�	��A1$�f��/o��S�F���sٱO��#������Xj�UyREՃ�`镝��ߡד"�S��"��%��τM���S��	�!,�G�4�]�,��l���ً��@��!�t�/&}fߠ�#䙎�3��\��h�^����T	��ۆ6�G$��e�1�gQ"�~�U:��2c�M�J~��g���\��|��"2eF�0N���E�o�m�r:��J�{$���_	�īu= I�O���`��Չ�.�4�8)c#j�i�U;�<��BW����E��,
�9�$�j� �C��'q�$qNK쫸�F�=�	�ζM�?<��hr0��4�:�J�m�n�� R�+AFJ�n�ԃ�A;��E=Q�-/w�楇S��K��$WO|�J���Nc��0u��N �}�������s�{ӚӍ�ݰ�U|�2�7���^�cN������z�`kR�Ɇ��n��|����%@�������=��=-d7���	6�Z��x�Y�}/uV�T�܄�6�	2�Z��H��K�:�u�w�=��ǅI����$s�7ԿJ��6���s=�R�T�[�v���h|�C��A�+�*O��&C,�OX��lF`Z���w�+{V<��!�����H�dmSϬ�X�͜wxœ�U��bݺOT��nW�OǑ�U�wnsT:@�3��
�'�iجkXY��K�)�2��[����K�͖�9(��d[n��ҏz���d�`(�1��alK3��*"��C����>V!/s��|�x�c�
�~�m��B�j&���z�g[5�zn�nDF!˚W�Q@:(�����,���~�_Y�%�n�O��!�V�W�����^
��G,������b�P$����B;a]s�����6|��w.��q��xWb�����Ð�%�ê]�H�s Ō	��;�4�����F�7��ZRSԊQ��%�Fc S2�9TKҿ��bD�ibN���;���!�O�ɦ��v�K0�є�L DX��Iƛ$��p,�]��H�g�X[��r�P0v�˶I}����]V� �^De��`>z����'��>��>�d�vx�$�0�hb�bᘥ򁳿)t�&�!��X��g����L�(?R]W�� lb����,�l��pI��>����t�	a��]9� ��F�ʠX^P̟�sf�C�E��@9��9CcZ�S��Kܛ��\�z��������fH�=�@�`��|��.��ẵ9b�pG9E�Ș��d7��Q��L���鏋P�<�-��Z#��n��i����(I��6���K��7&b/�pj�T=4���/0F �wq�����h�{���i�g�Gw����hI���]����?@5��y��Ʃ�I/uI���Z�H�m���B���[V������HG�A�,�a�d^#D�L]b�Ϥ	+(�C·,L�\��� ��l�f� lf�,���:�l��(I��A$H�	�TC0����<|���Ë���K��xe�_h�;:��R@����Q��J��T;����:���4����x�X�I;���\�}J:�Ms1(<S��k6nt� ���<}ܩ�ER^ׇ#���ŗ[�ŷ���6a�\���y�Ú��hB�0*:���r�tYQ���&�2���U�Q�����W����Z����I�ny��1�����>��j�
����N㠳97�?Q���AB���=�i�"�� ��QDM&����h���xjM�"0��&��o:G�����e"�� @�ɠ���k>������p�	T�s�/��;ա��݇ܟh�j�hR�#��22���wh�����ȩN?�"�,?P{��h�E|��jo	L�Jsq8/�^����[����5�6�"-"�%��-�c�UW?��b7�a��t>}`��yv�O�0i�顦�����l�*���s(>�K��}���-,�7��w�}�/�&�iY>�=�u�Y���e�$�'�;x������0w �	g�{D�:,P&@
��@��~'7ky��X��f-���{�SvX���ß��Ꙙ��Z�ZP� �\3�zdX:���d���^�B��"�+`��U�l&������leo_CD�w�]�Y���hn���������E�&?x-��7�97�����J�|��+¦��Ip�9Ք��E�Ѳ	�+�*�y~U��82�dd��3�]{�t��{{t���rp!S�o����>��Y�	�u��oX(4�=�v
�2�Y��Ӆ2��7x>7�)��4���3�^�����F�B�wE{���������~:��E�Ht���{��0�{�u'�e;�b���ΰ��p;��x�K�4����~H�C�[�bocD��8����*��3��mԏ cu� �ف[YC�`�'&K��B�O�㯳#�¿oS���p�^����).�.E$<�?	�>|���j��$=�3�4{T��Xuhָ@}�>R�'�C��0�����d�[�L}ޤvr�c�B���
ӌ�#l�q�"�ۥ��t����z\T�S�ܝ8=��U�,�e�Z�(W���̑6ü�ю�+TZ��]� j��u
k�w�#�M"��ח��I�%��F��u�u����F��ۨ�A΅�����-��$�{}���
��с��s�p���'�WY�d#���.�1���{��_e�^��a@ǮB)��x�P�6J��~��#[Z���w����X�Ȁ�A�ȋ��J�ų������Ђʧ�=�τ��8_��%Hy��-_���ϊ�0Q݁."�^���"�h�s�g�{� ���E>Y[�Q�YO�Y���f�.�t@�c�*�=�̮�X�{S�pr��Ac��թ�����%����!����7�%�c��G��Sv�v��aȪi��o���f��|���;���KTxC8���������;3���#��}��#?މ���	��?���
�Y��f��(���:Z��+ex2�S`���DwA5�x�7�l��ߩ�������6�^�Ä�<pQ��bA|[8���[`F��ׅ�1u���	���EKة|���,l�|���=�ÚD'H����uML_~�.XL��#"H�=��\+�GG��N\��Z}�᠀�Q!�\�,6#��;mrE/J��ԁy�-Ҫ����K�9����Zڇ��^���zQdoi6yUq^��):�K�c��Yo�N���l��h�1ַ��m?|��qɯ�1��;u F;1�Um��$���<�9���<j����Ÿ80aVo�3w��m!�I� �ц�g7Q�T�=�a�:�Q�����ټ�C�x�m�_�ه���A�;G�S�2hͽ���	^��*lY��L5L������06(�:O��/���d/��0��{+��ϾR�b�s,��2f�������P�u�ܴb���p*�{jY�����b�覜���W�D
�o>��@� ��٬h./����+"����3���K�
���"5(������6��|��
���@�Yêa�`5ā5��k�묂��P�>w�D�Ag�<�DN���H��2��i�f�OY��C��Q�n���1D������)�j�����`���F��T\�.P����LȲ;m�:Ů\����=�3ګ�n����,�c9�W��w�`WN3���zz�\�(�(&_��89W��>K�Be��k��Q@�Oa:U+�%���`�'���lข�Û�N��+9nt�i]I�\��<%���iy��^�v���J�՝���
o�[�)��]����O_FA�촪��!����_bk6^5��`��aeEQG��$�����������	�zOB\�si�FbGw�`�;�0?�����)d�(�u�����[f�tt�Ú肬��^;�ۖ��QQ��+��[c��/�BJ��\G����U(=X&]�*�����zH�x�����q/E�?k%k�����vɰ��J3we|ݜ)�۪�|w˜��_�ay}���?�������/�A��
� ���Ch�KA�^�)�h��t������R̓^:��6:���~Jin�J��GC��<���o�	�a�E��րC�'��ﷆ@���&%���e��h=h�l�^��G�i~�6�LT[�UI��es���g�Q�.�bʏW�=dN:%2��=.�\N�!���d,]o�V�С�}�\�Ac���ω�wQo���5TɚTm�dR��I��%��^�1������W�rṇ������^"�,�Aw�Oe�B�_ɐu�5�E����r���BƜ�T�`ܱr���?]��}�b�&�����w�f�r�M��@t�O�+��ٰ
�?�fOq�G��Z��� ��7���ɴ2��C��zq3H۩���Ja�/gT��r;�|ڌ}�p�����q�(/��D�
��@&�ql|9lnIm�Y��9e���\dnZ��]���{���xd�rX��ٔ�;;���'vH>U�>$Xe�񓪈E
a�FW�����ϤQ�]����M��(5��:h��܃7n� �!\s�ee�%Y=)���Oģ0<��wt{�Y�6���-*��.�@����,����T���YW�`��j��U�����u Qϡ���KMJYu_���k�#�>����4�K�G5ފk/R��~�4�c����J�B�� up��n^{���C5�6�g�:�W꧓ j}S|����~DM�uf5d�oh%@�
�P�T�ߏ��.��J�d�y��ϫpXh�\N@�����Oe��Ռ=��B/��@���V�CEO7�=Ok\�M���ىh����3�������MA�J�����Ť�y�*�T�u.��o�?����O���}W펺#���N�V��	�A��)�%�1��&�玻a�H;y5
~��޵|�y��	͸�iV�k�0
��$�i��*�e�C�����E�C:Q�\�4k*%O���a��j-�3�NH�I�OzGG�@��oÑ�}�M�Y8gؚp~_����6-�f�Y8mQ��0�ePq�AykGx�k�w�GǬ�2��݁!�H ����r�����_�u<�������?��<@.�^��Нs�EF���M7��^���5JIc�wexiE�`���Ϥ��`����d�$�(H`l�\��у���c��!�߀t����}Ֆ�[a��t�*q�՛�	S�&������-�_�و�%0��/wz������㭣;R��O����7(¸�%v�V�8Ğ���?���\@
���f���A��7�l&
eC��~��.����Z�ՇJ�3Ԍл�a_j� �
t�9��+;��v�I�[�Rtw�6�H)\���(jaS�`���4�<\,��[xT���3w���\��4˗��Zt��h��G����'���eϊ�����+Rm��(^_���{���4x��tk�m ��ٛ1�R-��%&&~�v��N2��Xw(G����RZ��5G�N�C@ӊ���TW��'D��������H�ͽV
iCZ�zd>�� ���i 0i�dm�iF��5�����)j9��;ì�;%�3<�B8�,��>����~�[ǁ�$�z��B3�-�X��W�{�t�_*�C �+Br�E����K��F�4l�om�	{�Է�����Y��'���C�M�K��y���@ze�F�e#�Ad
x��Q���D>{�IЕ,�my4���U�]�t�W�p7�˥M��qRw�h%�O�׼'̓IO|եyd4�QMxq�ɶ:A�)�Kl0��]C�T����ݵ�U�z�`,�ʔ۫3Rw�^oZ��gf�	�	�!_0�Lѿ�w�9�5i�y�b�Rc��pt�?Hs��*��95�+Fw.����Z�z(�"o�ai�&�Ǿ��u�L<>tkzJ��^ᵉ�*I����9
��sk:�o/��(/�,�<� 9�����h������(����>jդC�H��r|��LjO����,��}<�
�!���r"v�Fb����	�p5�^(�Ko��ka�q&v������e�w�T���&�J��<j��ʍ6����F�C�NʃL܈3�7�w��8vSGr�6��Q��"P��zek{�0o|r��s$ ;�����g)\���<�p>��g}��6�l!h��/�H����cp�iK7#^��&m�Z-xB��C��\���g�B���D��loǂ���V*�|�UV�>Q+����o#�_O"��0Gg�y>���J������i��(���,�-�4�K2�2l�Ꮭy���Yn�=�z%�:6����[�JC���^J|X������wh0(-�	$��S���߆���<�)u_:���f�	s�pg��c��|?�9�S�vZ�5�]��_�Y@���ִ@-���gq�e�3�&�����w� ~M�|�"����~�7Ɵ[S)�!Zi.d��Pp�S1��#u���漄�~���3��1������2��Dy6%�������{��ʻ`��x���:ձhƚ�	s�.��@�Ԛ9���AK�w�=%�>{�x��7g/E�4:�f���`�[m/����lEG�*��&�"���e\�@���/���g�TS�AZ����ˆ� �ue��
�T�5hW���#�h�3V�*�o���A+�b��ɞ�����n��^��������Fۈ�ƙ<���l�xa�ǝ[��G�B�@�2�;���8l����Ƣ�#�i� *���*�g{XQ�l��6��b���s#gގ�뮂)P�<w.�4 �U�U!EW���V��h|�FJ�;V�:�\�i�t�`�� �Kq6�kU=��C��.Z� H�T�9@�ȋE�qJh�'���y+���'�s��#��Ƀ����}�/��!El~�Wj�r�UQY�1�_Ш�mQ��r�Ap.2)�����W�D��<k�v���Z�����ظ��W��B�ȑm�,�c��+y 3|�2�Y��5`4�r��s(Wi��M1�׮�}g��7�~3OjU�T.U$M��Gao�#k�"���4�g�j�e3*lM(�o��-�l<�S��D����H�������7�������Al�۾`�]��~_������H����gӖ���	,�p�cQ�X�E���-�G�Ie�c���� ���z�b
��u:������*�3f-G�������%�R �Uʌ"E�<G'.���Ls\�t-t�VM\X�k'M�T�Ͽ0�D�)jʐ�:hi��x��ŋUZ%��/��`�['�D���,�(�j�&��}�u�/t�������t?k�J�e[���z��'~*J~�L!�
��2@��)���Xx���p�c��;��G0*��gտ� ����w�_o�>^�+���KJ5E�*��P�s�x]O�~���)Ƹ��-pٵ��rk S*6� ��Ofu[\#�r��ϵ�)���q孋N�[��j�(�w0��h���	��7�J5V� �W�vxn
<�����S��PTF���n�����h�(Ӭ�,�J}5/:�҆�{��(�4����Nb��P�TfԘ�LUv�ʩ@�H�v�3�&��T\�y2Q�D��;^b|H/wP#����P	��7ZL�8dXG�1D(b��ݚ'��'���,��7P՜on��Thn"�'�劰%�e�
*�N�;��X<�Ϝ�+C�N��8�ި���-qq"�3�zSL��V��
�* op���ȏ�s�MIa��S2!�h�@�u0@����9Ɠ��c�Ra( �7��[�y	���+�%�G���������ef���ˀo�{�h����^�6/:6)zA�z���֋�w��p4Ϋ���p��s&w_��{5���@,�T��F��.��,f�������e�9��ɇ�r% /UT����H�p�=�dO���E�}@Q+^o}/�}am�������3�*�CFq��*�Q�\x("�&��$u�5A,�ǕO��a�7��߀�)�`id�9(��e���_�f*`%�*sG��}�D��Av����<K��+&�� �%̣6vp`E��!����J�I�,΄��e�L�(9��be�w���i�&!���u�U����f��-�	�yo])7"�o�t`�8�-r�|m�o���%��qT��j ���QnHY�g�HRE�Bg\	�ހ`a
2V����=�F�t� ���sшS�{6EH�5
�;Rp��8����.�΃P��R�z�Ť 1�_���tMǀS�:���*���aL��|���!�<���i��/=;J'�P���rE��׿�/�;~
)
�I��A*�,3N�=�\� اB0�'�;�+�$��D��ԝ�ez��yͩ3��Pd|��L�dve�A��])���� �1o�nđ��X<J�5�B���R�hmj�)ækPd�# ��V�vm���ݰ�~��Ub&��	F�lsӬ=e!t�U���2|U���Y?�U|�e�>A�������4n���ߢ�T��������c!�S� h�BJ>PB��z6m ���	 ]�qL��<8I9C/����-w��xрx;�umF��p`�v�z����FM1�� ����<o��� V��_��| Q"�1����;�M�&8x�w��B�vd�}�/� ��-Aw����L���g1��s�=M��ɉ��N$�Ob�G[V��C�`z{���V���:8����z"�`����U5��ciC�TE��!ѥn9u]{���݈U�?5��rIe�T)+� �7�D�l{NTPn�Jr]��p�KȦX`�-k
��y�f��K��z���j�C>4�N��Y�Ύ �R6�AA'([�n�.��`]ޥ�a����)��[t{:�7`�=)wVz+>��Ⱥ9��z�������a��#���i��K�;�؀�mF's��(��Λ�!�<��3R-ҋ���EmO� �EQ�N�C�]]u���t�Q��N ?˃�u���N�nD��L�n;^��Ս.�����7 ���%`�:ż�ŷ���'�25�o8�yU���θ�%_ƺP/':Nx�V]���D`�g�&���#&o9ӥ�)���/H86��ς�8��0Ћ��ޔHEv�}J9��!T��)�U0�����0g���&�I�{�Ѻ�&)RD������UeC���͟�S��]�O�N�gW�0���Y񍬴�_JgXD�Ê�`/e�	�)��h�$h:z��i��^��F�:�x*و�|���#-f�̖��� �������DY`Wb����1��߀(��Q���4/-P����j�5x3`����r���L�8a��m�gGqs�;o�sf#J3��!��>C���P���ڕ���P�}��.�Ze��k�AM\x0�ú>/�t{��V�q-���@�Ca�t�|'�+A�>�h5�3SpdINv�؎a��������u������i�>�
g�ӄ��%�w���3s!���?��}�^ %���=�md�@���[_��Q���O��d�*G�n|�$���k>3���V8��^�o���>����I�����}��ƪé��=tޜ\
�� ,�Ǒ���+W,���_�b/ �x6�mV�j*@EW�@`��:Vl_I����EױE��ۜq�GRt!XM���ba�iUJGO�SX���J�
�k9Q��S�ym\�x���D� �q (��{0~��cz��s��o�Gx�Ƃ'A�3��9��?(j^�n-�w�h)��5Z��xs�Xg)�I��R�]���\̮^����B���)��O��n��-3�{#ד�&ي����4�~��[�>5	�_9�%����&��
��D��E�j�Y��H���aipo`Gʉ�yf��)��*$N��H6���O�X��/d��E�	�9��V��)��b4����g�^�����n�=�b�Qk�꼃J�G��+�@������_�p���!;�)nV=�r]�G��L���/0�?Xz����̎�h� W�X}�y1�_�_����m�C�b���n1�.N�"4U*��ц]�k�EOH��t��(��_��B���N���;
�?�E~�o�k�o<6�]�Sw>���ι����u4CVi� ����[��EEG�)	���ރ�84�ѽvÊ��3$Ƥ�!���r�Zw�W'�� b�H�^�l-K>���u�ML��YS�p_?�C�qƑ�^8mi�'o�DJ���ly-"cS����u��{� �	z#[�e�^�� 4�,5��h�o
k�Fj\b�J���1vڹ���a�S�H�c���)X�'�p~�#�Jz���Y���A�"��ǹ�mJ�� P���6E}��~�������-H�O㸭p��D�*}���佲0_u�q��H�����[������=��p�)�\,E?y�>��e;�U(,��#� ��i�4���'�����B�|BCY9� ��q�B��͈������31;�W�P/Xj�N̘���I�tt����	I-�������e��K�>��C��h+���(�}jd�P�x����GL�e9�1���Y�4�'�����@�.���$:U�ȳ��r�)�4��j�~��)ԥ�v��X����E���a�Z�P�.���`D��}�G�$w[`a�%7�<n�R?�M�1��Z�Hm�,٪ ��v���5S�Ƙ�0�+_��N
@�e�A��J�`�8��PTZfS���\i��'�VG�;B���S���ʘCQ�d�~,� d�k���:%�<'�nE �p~�� ���^xI͐�:lTDЙy�8X]p`r��t���&(p�f���Mb/�N,EH�d��&؂a����1
]�i��2�!:H�:��{���u����u;��zJi��5��4~%5��J�gv4"�-�����&6��9�E��'��<����=�0�ȽƮ6|�nN���X���3��i�G��Xc�0��>��m�GG����%��0����w��m
�������ZAh}.|��B�����mm*��vT�vH���8��R#	�NS�^ϙ�-v�ʰM�<��-�x_��=�e43Т�	R�%w�HЃ*��i@y�Ecݐ/ﮏ�e��#I�5�uI�o2A&}]a��'0K�Jk�V���h�+����Z�`�o!�"į�L��������f��$i��)�[3�����J�?mD\���UQ*dUmk��kN�5�ɷ6ʖ��0���#�n���r�^�q>F`���'J�Zs	pFy��nB��~����	}���d� 	7�)%6	9�� :s��[���U���a�G<"z�DG�t����w�
c�p�4�dL�*)nk�M��k��UD�v���׀f���� ���|�Q��)	���Ơk޻�+��*k
	b��5��ȩ=��!�)X9�PX5�D�,O�\D�7���ä9��y��9�VǱ�J��kK0�C��;HK7P��|;��dq���G��g'�#'�2Vv�.����K'ᆝ�B�SXR,����?q��|u�8Y��R�ʤzѼd�"�
�y�c<�K3)�� *Y�µ��޼RZy�ŵf���LҋK��"�]Jh�'����7_-l+��.\.m�vI <?�����&�!������~��&��A��Kx�W��hE�V���B��uh�U�a�)@��	9u�G��m4�f&�ߗ��ncC�~����Ѽ:O����|�1�TZ=�O8�?��0�tIc�ޫ��w���zg��H����B�x�(�'�x��*�|�y�E��gQ�SЭ�3�ɳ��w+��ӆ�lZ�Ю��vzZ��:\^��M�̺�򐉝�z������{�$��/���8'@��}���4����`]��$ȑh�s��/D}IX�\�h%U����Qo�78U٧P�E�.�����p~Z��y�5ɚɸ�$�����i��,�&��"\���\�u/����
E�nc@�r#tVr���H(I9�;a�g|�'pU6m#�k�s՟>? C�|��	��E��˺7�?7�35`�*����.48��|����}v�B�4½q�Ԛ�/X2ԙ����U)Hw�i/�]�NA]�ٻ��IK׊�1��v��ߘ#sÿw'{uR���x;���J���Zxd��d$�\�1z�Ԇ:_��=g�'Aq1�?^:qJNIH|�[�Ɍhه�����,�Z���yc�iO"cf@�h�*xd�r��u	<�K��\������|���l��"�1	o�/�P���[�-��*��e���7�4�Uǩv'�jC�	F%Zv~� �����H7�
�"	Gݝ�Ký��&���'Y�4V���6�Y@CΦ� V1zȯB��H?	M�OvԾ�x��l���g�&f~N�G���h�f�0Db��1���
"I��g�r􁵬O��vɐC��`2����nB!�`�}�8�)��FXr���J)���V�gz�b���W���B���T�p�������>�ծ(]�!�>�s��`��"�7���k�|�X�'`�7H���,�	p3��M\F@� �.+az�h	ۂrD��s�:���@��:��j��\�Tp8��rՆo�i�k����FS�cy*��:	�w_�a'���1?c�5G�G��<�=T���������(E����M �2�ԡ�b겄�'��L�"��gy�|Ӗ�5��sG�ݛr*�������U�����L�br���s�'p��iײp)���~��hSi,AƆOE�%����a�.��ڢrАǜ'�n�W�UŴ�dA��w�z��giP�V����>K��[_�i�����IU��	8���e����BQ��dU=CR��]�1X�q��p���cq;�P�ߤJ?f4'SnI!�f�U�ľ#���D!`�>���s�,�0Žq����ܾ$����
~�3�~e��ע�����H�zd;>�!�;+ɮ|��iFN���[��}�leAZ1�=!�u��V���:�8����d!��
���u�wA�Ȫ�3��u�/��e���)"�%�gS�a- )Rq���G0�ާ�UA�<��ƥ��ƶq�WǗ�-��߲����V�P�;���H�m���Ib�s�L�Ύ$
v��7q�ݫ���)��1��$��G����
��0Rg�=�f�۸��g�Y��l~��%���
7䵖c��ǚ �,?�/�M$R�p)�
z<[8,t��"����V��b�Y 	�8����&�>G|���5V����:t2f��O-t�ꖍu��d*�XN]����2T3d�)d@^W	�w���f��v��K��]V�A��ݲ���D��%�.��¿Ĭ����N8o�Nɸ �n������y�z��<�5ҿ���K2���9�lwnky�Z�&~2�7��j��kT��`��? ��H�&iAo>�%gk��c,??�JѲ�y�i��>�b$ܪ�p;�R�$���s�����u���{wwC��#�e:��y��k3v����t��!?�u�q���r/짡�u#������&�%����~�1o������Dր#w��M$�@������.zy���� i�Q�;�މ����������H������%�ѥ:�4D_z����m�#��� |>ah3���.�fY�]���'i��P�#g'��������(W�¼�g*	�A|!c����B������f�H��4�m\e�l��q*_NSؚ�q_������DPP$萾���Ǟ���/�q�8����}E������+.t,Fb^�c�-�#�L��*uA��ӧ1��<��'%�*����Uq~ŖMxNO�<�{$1���C.l���I.D��P.��ch���"�ߞmHTKg���!��F��Ë́���Y����\z��b�C� y�3��gG;�?��i�]�7�a���L�!�w�8t�k����y��4\� �*�g<�-��f<ڀ##��h�uW(VS��x�����CB3we{�.�t���	��Rc�L״���U?a-�dY�̏0l��
&����穵��K7[Ɲ��*F�x^�S?NF�:���gMNeU8��{�&�B�'�.6tǟ�}�2Z�5țjUJڝ���>$#�>�$b��:�F��8���p ����ċ�A�i��^w۰K�}��Z���E��{��zx�\���|L=QZ��2�'@���v�v��Ǥ^Uz�es�P�8c��k{� #+�!dZ#f)A����c8�`�:��E~�{�{��b	�@Z�,G� �����"C�6�5�]�߉��JŨe�()��K�ʵ��M�J<.�3X�Ċxu�ZLb��Xm���Q���7|��h�Y�z�b�j�CG�ѭI�m��a	�Y�c��+Z��KM��꾧!L'ߤ~�Kݙ�9\���񬢄C���4�b�+����8�#� ��	@�ԏ���H���hS��z2��~U����E���]1=�����bɬ%��%	�0":?�>�1�� �U��l���Ɲ�CL5��l����(&����2I���pL�	K�n��w=�a?*-5f�m�X��1Zf�����#_�-o:��쮅�P�zٞa4��/DK�X``���5����hBZ�ɦ��=v���J@2�\l�[�k��WI5+��D
ra+d�ga�<��k�lg���-���Ź�Y:�I��_��Ҧ�I�
W��A�':��J��}G�+�7y��]L�+�r��OM� ��-)�8�Տ�2Txs��q5O�v,���~8�BPh0�����ZH*5�r o1����|l��M�����*G��#�]�wT#7c͙K.(r��=ʜ��=1�I��gIӴ�����d_v
��0������1(��x�^�����@���9��b�����͓�|?z����O\6��H���;ȁ~UF�7'��]���T���V{QI�>���:�y�����T�C*�_(�mt!ϽK�:���:�^&����K�%�T_�[Gg��H����+��������}��:��������~�[>�k�i2���sj �~����y	ڔD�ęMV?Rؼ��W�֤�lG���Ҳ��� �0�#ċ;1�����x-A4Yh������V��s2o�������:���rD��෋�'� ]`�o������/xC��&��?�W��r���$��we�����xAQ��$���K'S�(LV�u�%�G�ސ�N��@ik,�S�%bNa�����z3���j�'%U�g"X����"�K/K/h}(��q�;-]+ܘä�����ۗy�X	�j�1Y��=�/���Ɔ1}�E��N>��/t�q���OQ�U����J�&�B�!��5#8ZKP礉,@���`�-�49+�8}Zp^իtGh�^w�l۹�܁.�����-[�l�Y:��q��%:��DG'Y+V��#�]�����F� �w��[��m�\�o��F��y���O�iכ�o���r@���%���<Pu�	;g�0�g����g�������˝O4@�cc�-i �6�_)��x�ٛ���	�1�p�DŲl#�:�����gWg/O�c���� My�t!!����t�{/,��Y�@�hi�,M�(Ǧ�{C��F;~9������gu�ɕ��'c!�A�\K�֧>��@R��%sc�~��Q8m�7����g��j�^j\�&�7��!��!�9����Z���3�/�A��8,��F��Sy�g ��C$Ku�0Y{ôB�,�}��@7���:��1�Wm��执� 4��^ni���>֓�ܢ=���9��5<�y|������ֶ���Q<��sǵn������N��U�����R�V��(͇�Z����ï焵���{��4���vr¦*L��9G#�j����1�����9���n�e�Y������<+D#��9 �|z8S6ΛB�W��Z㎳��#�����������f
!?�A7O��[�P���|��݈�ˠ��ƚ����\�u���"͓$��8���㪇kv�͑9�߈��)��ZAdz�m���q`NO�!���>��^'�g*�.�X��vv����K��l�2��%�<k����
�����G�&X7��.�bI�@j��x��=� �?H͓Z�'�9LԈ7�rw�k�����?	�~w���Ŕa`3`��cn� 2��~�����Ka�̄n�G�|��������3��<L��� ���K?¨t�� -�'b<�3jp4�֝O�nT8�W�5	���nF��GiH�'���G�Fr!�rӕzf7^�2��s�ό'���U���n���7��<��M(:ۮ�����W�,Ht��ͼ[��t�΍%��!��)7�����6�%d�+ӗa�(_�[jf��*�$On+�$�x�g58��f���W���2��0�r���-�q��>��_\�hJ�`<����Υ-Q��>BT7�2��y
8"�rc�ݟ�׬�i/�-�Mb�/��o���/�r�����@�-�Z�,U�?��3�.5^�Q�V<�33*�O�E`#�2��i��e2�ku��ۣ�b��)�0����q����=^�}��$c�4"�} ����a]ZL����q`��K�ȅ��l�̑>R�1��Ԥq+�� Fb���;,z:,+��_�@q�a_H�����n���m���G�ޙ�����c	D����k�]��3���	�6g��T��zSD��"Ln�)RW\�q���5��ewĞx7��98�rh�ܷ3�2�4KiB&��I��{BN�L�Z���8K(Bb  ����f}4@�#t�t�QT��-�%�'e�Q���ZA�R�����9 O����0ɴ�,U;�����i���f�䐺?��QB��S��O0B�iue�hW.m���)��E��o��=)�h~��nI����>���!�ܩ��;=��]7�<c��lS��� l�`��*���ΈY��)^��nk?����0|'<2�&z'Xm��ݍ����\�q =(�D�M�{͸	#��3?�V{����gֿ����fj����"���p ?<��re[?t������+��s�aq*��>zܩꎢ�����D+.Lnj�\��oZ_���A`?tA:�(p�ec5z�*��n�')F]3���ޢa���"��uow2�;��<��C�#�s�/�m
_���P^f�����߸ �����i�WB�yGϝ����������C��m<{�27ȅh�[4C4誑 �4���b��U:���!#F�ɺ$y�8�$�_;��;P~�ɬ�e�TU�n·ʖ2�Ӹ�Q�i3�@� ���R��҂���]�rd��|�*͝A~ڕi���KQ�v�՘�$���	6������9o9��O3�MmJ~�k������Wc�Vn;0K��YMP����á�Q=9|�?��i��@��¢6\n��g
�\�#/n6ʰ�Z��F�_�͌��j�:�k	���cM��7�k�O��*�}jmc��W�ӈ�t��[%0w\m� ��asNq��_�Y��N�?lu
�m���bH�:��q"P<�����+lg��]��
�Эt������"%�×.��9�0g�J��;�b�t5#�dy���X�72� n���O:��Lٌ���d�����Ț�Z�����2I<��UCP_���ƳzO2�o�H�h� v;p��}k�c�ȕ�ýh�J��A؍�S4X̊�;_&P���4�{<���[C�㍇�'� ם�)L#���w�`�7N��Fi2?|t�y8W��	�Y�S �������/�� �ߥ.�AY�����,l�R���R�/#�o��K�|ڠ�����6ʅW�_S'/D�y��t>�\��e8Q��K4C���>+�rdsW�P�Z
tWzPݟm���c���B8g�>��%ҭ�O�(���u����銚�B�?���+���ܯ�֧T���:z�Ε��3�ڎY//���V@�͞��*����>7�,���U����Y�̒U��)Ǹy*9aL.��w	`�q��u}{?D:����<�vA�6��?���"k(�_3�mTY͕��=	`.zi������0ٟި,�r[\x)���a��U�2	st;�QbK
H�יּ��D���Z��i8��6A�ʄ��#N^�{����Ci�;�8R�I�U&dW������On|Qv��yR-0~Xgk�v9Gq�<AL�|վHz�y�A-��Uw�e���>;z�����)gCVR�͎dhwF�� ��q����3>,�#�kd9�̞s�Զ5uvU���kfMƆ�ܥ�@��{D��/���i�d�85(���#���&lNN�v�d����n7�x�� �u��wz3/3���)������"�b�ɫ��	 .��O�6x䋯�]����eV��с�0;1�-+h����&oVZ�r5@�#{2����܂��,[��l����(�?6l�௯MD�_t�RGtņ̇T�����i�N0���Խ�4��|���צ4�X��˫}��zM��m���үh�X̆D�ЈNΝh���s30B�1LE �sP�NuT�q$-�u�_��>����6��$-���{@z\��SɖJn���g�$���n�U�'9ě�{������(�XSk�Ċ��h�~7',���5zx�ٸ�m�����]5�,��8GQM��j@�^{�
J	ĆCN�T�Ra�b��=mU��0:�oQ2�Rf^wa�C< �G��^����-��د=V�!�q�e�	��&���E!�WI��RoV�����L�m@_y�b�u{��Du�mk^�|����@&��Oۣ��c�RxC�~B�8��l�W- 6
{$~l�[�.֍�j�lK����I�Sƚ�j?sK1Wv��H��<�˯Nbj��*�ʹ�� b6��hgR������%��X��N�#���ꖆ�Up&H����{�H�Ԫ$��~�E,������Q�X���l,\�:�3��?�p��8B�Ț��!v�eFW�$j��D*6y'pXj77��KcX�.�ɚ��nJIb&�f�����u�Mݏ��<>�$��F��i�D8�N���Ҧ_2��˿B0"�j��eS�4)�CO��X�j9��'��|�jv�7M夲��j�I���Q&fx��A�m�QZf�F-���%��V������t$b6��U��3�m��j��t>��mӈɝN���X�l��w$�����[�삒���[�`��CP�Q8FBQ8�����9�{�Gˌ58 XS���c�*�Fݏd��W#�Q����6����p�{P�_�b�d��16A��\��4��^ϊҟt>�$�j]�����[~M�IǕ�Q�I3�6YNv���&����@���(Ѷ�b��
���+u�Sw����f+O�ڔ-h���p�+��:+�b���,���s��8r�(��}��_q�������4�L�q�MǕ�O;z��y��`o	($��+*�順���.��t��ɞS]���a��e��0?١�}m4�1�`�󎅵;u1�-� ɂ<}ਲ਼�>gL/q */�2\A�� ��-��%��5Aޅ+��J1�H"���V�����g�N���*�=�'G�����:.,4짜C8���*���	L��J��z�����i�+i��#%�m�,G��5sm(e|v�j�%�V�E+"wf����W�$>o8��\wrN-�^_�p�^)g�g�?�	�LԤ�"�OokH��B[����L�lvÊ�p����ZKˡ9,H3l��^�}=�x�����>�|UjҚ"��Ϲ��@�UY�٠�jͭ��Fzn�P�r�n�q���?���,IX�m���đ�ȦZ�P�|�~�]�.Z�
��g&U�0�,���\�9η�'�A��]%)(f�W�o�����%�A�ŋ��Ù`��x�t^U�h�QM��N�ox���h�9Q!/��ڴC2��l�.j�.!�7�<�c�����뻦[Y�l	mƤy<��������
�z"�Uf�Y��H,S�CP	�zĖ'0#��|�E�bچ"���4���VC�Mr$% ����d(�E_V�_���fT�`%F_5�f�t���*��^���z��nLB	s(�E ��J3i�2pa����؍q��~}a�?].I�^.N���N){Z(0�!/cE���onqxC���3��8ㆲ����~%t�\n���;2��v�4���`�Fz�?�؎�уM.����k,΢{#�ߏZ�_o�f�5��oiQ*��ԉ%�sd=��G�2A���?2j�������v*SDI�G�.�!�U�+�]���l/A�x�"���ހI����
�N���g)�mn�����0ֈ�d�?� N��S����0D��u=��ɻ��׎x��+��{��<%����l�k ޛ�Uz?�{���Ɵ|ע�[c7V�͉�U�j��IM���-����OB�F�G%����pa���/�:/+3w��i���d���\{�Fx6ͽi�R���5D�t}��ɩ��C�IT	ͼ������m��S7�Mh<-|��~h��Z����!T�[(l��\Fe|w�K[���.L���+�ճX��hz_�y�B_�b�����6�}m�B�[��Zd,��+�&��O�*7�~b|��?C����AWN��v�FA�)����9��T���|��~�4�[9��<�Y���'_��?��#�k���i�0x`��{�w�lʗ~Qb���*��y@����&��F�-������dq*��f��%�v�&��Ph[%��A���6�����SX�L|OT����Z
�{|ܢ&szw���Q[;�U�DC�D�4�����U�ޚM��=UX�d��i��݁-Z�x=&Lس�������wsSq_�S�:N�������Q��,Rn`	�;�W�F�Gzxm�2(M_X�}|;뉆d�ގz�+��U�&�`��-�b�`O穚q�N�4�T$����i�.�z2��m����d�=s�s��,´?��o�K������!dE/��z*�m}�WjH�K]S��~�%L���
]zY�|"2?��Xd]m��O%��m��ѯs�t-;b$��%�wu����������࡞�4 
�f�<۰��~'$��MH�Z�����G�Z��Q"��m͙�d�1~j��ŝ_.q0E�ʩ�`"b�ܫ��5�i��:�oF�̾�ˬ 9ա���V��Ҫ!/��0�5���Jڲ6e�J�Xw�?l�Ԃ�$�w�r��p��u���w�ߟ3��.�^�O�gq���3�| M\4�c}J9�7�~&���� �����73[�%��&u'��׿�Zo�1l���#�����㽅�=A�G��s������s�hn�O��z��z��V��3ti]S&���2)����y�T��}IU@��v`��1��N�4��T��LǦڱ�Um��P��V\[_k\5�$���zv&y��y�Oɘ7*A��nݼ�?�ɼ�pDD<FXs��UJA~�`b{:d���<�q���y0���3D¸��S�>]���!��^�5���[�R���ne����jg��܌����vS|��z��u!�.,��DPq�@���㺠i����~i��i�� �N��_U�oac��BO����E��]*W~��S��<�.wuǁ�Y�����M�k|k ����y99�K��f؄s�7�8�ͯ���t@4h	�2"5z�k"�x�&�5���^�x�;�^���3���Ժ=�J=^���T'>�Dzɔ�����L�3��˝�	o �L�Ddj��U�h�M��SnB��B���[�}KAփtO���]z�0�,w�F/�n���J׷����pg�v"���Y=r�Q�O|m�qwG�Wv0��I���]���f$8�*�Ĩ�H?1e2�k$$bh���ٵW��ԡ���^�9Mx��qR��6~�� ����g�c�I�׵�z9x0Y�d�k~ތ�ÔZJ�$ن#i�OG]v�s��k�"θI�!�MT*26e7�j]l��lC�p8�'fY�%�k睰��F���ίV|�䎎_��b_�|�p���Ɍ���#�~�g��ܥ��Ӭ�mh�����}s.v����"\2R6�Mv�I~5�-�o[�]P��U��q޾���e���^g.���?��w1ԓK��lJ��D���a��{Q�y���^e#c����<Ā��E���}d��"��u�� �%����`tuN��T��" 3��+���h�\�^ �e��AT���g��o���ѩQ�5���ÝH�����e�����B/din����M�,7��6��&(�X�^t���/�m�h`C���ͱ>�܍y�����f�d��oi��-�[�Hk��-	�m�'!/z�
~"+Z�}Z%a� hP!$CT�͔����"�����1]^e�
�ZO��{W�s���j�?�_r�P�<� `�i�W/�2�&�3;�<���y�O��=�n��@w�OtdQ�H�ߩ�gҰ�Ȫ�p�z��6˾
��W��ʾZ�ʒ!M���V�j�x"���ܖ@8��:Bh�;���l��C�[nŶ�&�1Sp���!��;mu^�'�}a��6�}���nt�����H���ݿ�H��b��8q����/?/�*�ơ.zP�T�Db~H�]q���h���Rz��� ����I �x6�ǚ*�@D��EI���6�ҽ��[�QL����:�}��{�^�g��!��1	QAؓAL�@���E��4?B�x?äp0�/є\!�&"���yhYW����`M@��R�h�r̋Q9��|�Ŝ�c70I��m���@u�@*#�/���sR�a�yU��W-�/T��7M��7������ۊ����J��Ȝ�����$� ';�0�L&�@�u�ޕ쪞���J�feŃmT^&O��4�r��>!o����r�޸��u}zFT�xt�SՐ*�e�lkY�a���Vp&;����v'����]F~�9����\b� e�(�p�w��s�����HA`q(��QJ�E �mg��r��	Y�)^ӻjk����]	�y��/
��~.��Sy��l��f��Bz��,_����,蘢<�V�8�������K���!K���8a�a�c^�L>��`47Q�f����8n��=z�N���|G�?td���@���,�jy���$K��'(�]ݾJ;K-Z�1V)�����	E;��ub"�_�~Y�p�	�����ՀDq&�!&��v(85x)��-Opύ�� �dL޽N#$�7��,�w���df:��n�$Q�GURz>�����E���|<�ƈi!{�q,&	Y0����,Fǣ�;4#�SF<���^�k���Q�mҘ����> ��Z_�x�\쩵��$���w�(���s�S�7�X�cL�qJv�|�H��r�ל�2O�>ivk�s�Hڀ�k�2�
Oz3�5�6�EX'9���u�a�� JE�g�'�0���bh��gyQc�kؚ��oc���j��A�T���a?ҹI���������X�>�@/t!r3U������ilG�kɔy�����9�XZ�}p�XK��� �0!��rn���yr� �6k"�Z�=�a48|kkZ �E��P���|b@��	%1;�����[	8r�4
���2���L�[3O�j&��k����QnώVr���{V�$��E�3�P9
��Q�n���T�reI��Om��34�~gx�5���ƼN\�IǕ^fF�g�N�(ak��~o�e��_�`Y�(��-��!�8�Ot�d5`��l-"���@��	�!z#��3@�P��(��+�@���1�؉�M���x���ք2@ ���z7�S�_흥R�}	?Ik5�#���&^�U����	�u%�V]�C?l�N�F��ǸN����Ŋ���D*��S �Q�1c$�;G��-�lR��n�[;^�n�:���!��h����{]�݈GO���ex�yMbG�F����
�	]�dP��?�R��iOX�/�R�hd��DL�a�k⿓H�魸��UP����eK+�&u<�FJlM�k��GP�cg�EW,��o��%(wW���V�L��ł�{2F吊6�w�S`B/7x��>��6'Ғ3��Ъ���V�Z2��u�K;��E�m1�a%ɬ�a�gt&����ܝ�v��il�	����|3'���Ks� �x��sh��wJ�
��"^eH�n���
�񢊹ՠ
Ip3ߡZ��}���L�K�h�Aå��JM_�"�Xߍi؏�]}�Ʌ�H���w;�9ʩ6d}}�)1*�8�	j'$�2Y0t8ev8/���)�j\^��/c�i1��� z%-� �e�.U��r�[<x�"�ն��������1���y��;Y\�7��f�)��)�9�@7�2ml�����9���e�x��� bBA���\CA��ы����c)+D�ʅ�!W��(�\I�R�y�yz�������G0�
���RY]*u�drZ�vU��9I�G�{]�cۢw�Ӭ܉�u�?�މk�&��� =�-"թ6�ܩ@�P�u�{��G���3��]���� q �kT꜐=#������Gϥ}ۮ�CfnO����^v�6�]��1Xdp�����DMF������Twx�p��.����9�HG�+W���%7����(�'���x��g��ݔ�o�ys��D�/��;_g}J���۩��4Y�]FY�Dۿ�-�h �E���΀,1��}m�9榌�[;�M7^����մY@��#�?�k:]{Ὣn ��+���>IO��q����#&��,�bTJ[��Q��u�k3I�pyoS�c��K��\����R_^?7J��o	M$>w������3o�F)�]j��Ưx�,�zg����f��c�@ԿE���m��7����S!M�yZO{@�~ͥ"�w>���J!v�T��xѾ�/��O4n"�����N䒯W�'v{(@$0��Ҟ�{>j���"+�|�1�̤ �*Vm�:a�´G�ag{���BMbރhZ�[��w����J��q
����ϲ�}7�ce��]k)�}7��F~X�':�,3]�x5'��:�K}M����A�ƙ,�$��@944oΫ6d�hO'|�/�7�ˁ%��G0w�Z8� ��1�g�0p��  �1�@��E����
�~�@B2������k'��� .����Ū���Q��K,����9`��h9Tّ̏��'*$���5^|.ԇ?�-��w+Lx�DPY�͏A��v(��ZF��d�(S���C�1�~z�c�f��6���ݹY��ٔ���TK��d��]�6[�UO�kG�,10�>�L!�y  �Y���`?(�q|'|p�˛F����E�&���t-K0�q1>��!wa%\8�������.\��=���҅ZBIx'�6��e�o;*�n@�P��f�E�������s�^{�@e�9�u_�/��[m��dLZ�(�h�MX��	�[����H����t�a��.�q`ƂNB�P����3f�Y,G�����P9�9�Ϡ