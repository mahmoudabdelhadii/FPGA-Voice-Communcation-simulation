��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��,�y�}�ǰ�=4d�H���`I"��W�`r���T:tB�T4D�m�)�	1��I�t��
��8(�8t>s)ו�."[�漆���]�~�]��;�O(1#5�-� 偙O��QZ��~rL'�x[�i,mׇp���O�I43��4d�,�H�����SN��d���3���r��m���̨T�I;uj2Y� Er�*p�Q$Gm���p�V�`�2^���,hz�<p��l�Bxt�5��s��\yq���#�@W���f:m��T�	,*�񞭋����_��㧋l�	�\�:��uGd��PǷ��N�I��_����Tuv� ���us�(H�~�{2H�:Zor�Q	#%�3ˠ!��iS��95�,?�.���/�F�i{#���Tp5����Ҥ0{%���2vpn���X�����@l����3dc�ק�3	�Ed&3�ZN O���z��s�yxӡt��v*}ԫy nj#��lc��m戭k[��5)�A#�����8�!�]�Z�s�M���t��w�!��'ÒE�rv��Ϝ�c@<U��\tq+��&|�&X1)C�����r�A~��B�&�����s�:n{p��͠R�X⺂L^��R����c���f��J^?��ܣR�O 1�rV���:��T�4���AD����˩�F�w��)Dm�O�b,�a���1$��c��7t[i2>�ޔ0,S���󧇳Ϟ�ᒨ�-��}�!6��Jyv�醊�^_�(�H�(y^����o#����X��3-�k\8�M�T�"`R�DF6ȕ� �,5�;Ҭ C�k���1\������k�t־9�}���� ���QHF��"��t�9 ?��{E_�7��!����](�S��0�q��w�9��=�i]�1�GʦȪc�W�XC�|�$��}q�6����zf(�u�� ��lQ�m�x�`�)��O�^4ɏx{A�����i�sp~�[i�nN����� �?���M%O��[�-�: A�E�����Иɫ$��w�C��-��@m����Jx��u}�~��;$:z�����+�)pEH�@59ۜ�&�1"W�ںٛ���%Q�P�5�$�#����L���=��w
��ss��̔z��u� �ˍ�z����{���zZś�j]��#ĲwL:-������܋L�4�f\�v�fae�~�H���z(n:��Zn���{��	i�£ջ�/�+��� ���<��:�9���[c����F�+�v\M��Q�nD3�:y������k�T1w�tyF��~�,�ӬV׀�>�љ��m��Z����W��(�$�I���mD_�f~K`OUf�� �vlr[��{�[�8Tl%&�����(駙�eM�;^�.i~�8�����S�Ke8���G&�T�o-ۈs����*u����Ȣ�4��S�<����x)`Km"!�T�31�)�~�ݶ�s^4���@�Z�*`��̺ǂar:�JFv��Ȍ�|�K�H�'Z�QYy9\�8�K���uR0v�N��Q�x��g���v�p�\�!9�9�X�F� ���cX��ufR�O���ʲ0D�n
Ӷ�(�p�Y_�:�����VDf:���qA�a�� ���N�\M�8Y[a�OT=;��D��@];z-'������Y�SC":g�?��@_�+ʙ<��Q��V�`j��Ͷ�Mo���-�	$}{�2%��!�������l����\V
gW�i�T]�����đ|:!��x�Rp1��b�'���@�z����<z�"�e'��"^g����wl6���H��s �;���e�qm\���n�K�]��>̺��������'x��Xd������`��N��:��bX�:�	��.�S$'0&ذ�{�
�~O�X�R��.�+��ApX5eE�ڊ�E��� ��<�k6,��J���;CP<m�����ZRޓA�#*�,��=��K���t�(kI-��4���
�.{��c���.��Ϝo>WY�^�z���e�e��`�� ��7
�۲�pJS�����7���qª�)���epE����� )}�x K쀗��^��=�JG/�@�a�N�^A�j���ɥ%@{iۉ�Y4�Bʼ-��+���F��#L�M�
�Q�zl�T�댌0��T��%!���s��uLSk^&�ڔ?Ϊ�iR߀;D������\�/xG#�]9�F��O�;Z����cv�˱|7���D�L^5�~� ~3E)S��{O_�I8�륄�`@8���݃�����Dh��b�==A�}��:`�I��~1l��E��틙��9�t��;�Mn�P�$�#vH���5�P�����EБ*|�&�m}�R�#l��R���Sy��w���_Ӭ��p�06��k�)Q'�i�4�c�x6A>W�D��O�_ ���r���3��p��᤮nQ4����U��9yz��VI��@<�q��Ym�歈�4�a b��	 z���dh[ �'�1�� ���=j�������v�<��*#��-���U�4O�ٰ�&��te�ё��6,v��]<���yzM��%�])��������~򷪆�3��ey= A�ױ��V�� E}~�}�XW��@n�S?ӭ8=19�(�n��g�;��h��`
&ڍ���k�=�<65��ؒ����}��N��Ym��f�x�@uV��Z	�vZh���!��l�]���+��īI0�Cϙc�ډ�g�ԾH�o�:8?b���O"+��&���#���"d2�iJ���QA�-��8���؎�[�Ά�ܟ34'�a����1�8�T��Ĥ&;��n�m�y��I� �tq�#Yt�QZ��XI�J�L�G8v���R���6]����NFDmQ�:v�4��(?Ԋ��4g��Z�K:��d���ϠY�Z�ō��(e͌��Hgo�lr��Ѝub�(�-�/]�$|U �Zp���[n�O,�w#<�C�>����sgLc�m��%Z5��¼�4�a�����0�������SJ9vL.�}��Y���I@H�h���_h�#�s�Ӽ���P�n�6�Bl�Eġ�D�_�d~�o��Ss��ڋ�Fm�f٥���Y����)�ej��(��;iy&���|+��AQA��7��#../h �I��N�E��I�5(�����Z$ݣ���DW��/૯G%��b���,�TÅCXj��!C
:�b+�6޷C�Xڙ�%F�>�42�O$�aW;�����]1yB�<�5z�Ӿ̕�˓�6�\��+Bne�3�6t-˷�����3�a�l�l`B��Ks ��;'m�Q��g�˨A�Q�F�">m��K���jb|�Ҧd�R �Asµ�k�5�hu�w��cu�d�gߔs#�Ӷ��Rp�v"Թ��ݕEA�:' 6vfB�5O/m*�vS �7?!�b�A�G{��_��-�,��|���he����,��dǮr� �؉�������4��Uj��˞e
to�j����<u/���~�%���RSA����Vi���ګ�2E�q�i�Q	Mw1c��&�0�{�E�wmd3B5��m���%}�&�އ�<���|����(�L�u�Ɓ�Ǳ��ģ�k[o9��/���d���4u%���o\�|G�����
�����vI�)'�w�� ۓ�u�������J�'@}� .7/:�ȁኡ�E(E�q�zIM-�����r�sRe�K�<�c��L܍%F.�n./������'˶�kt��jj�|����C,�6�nL&���҂o��Qi�9hB���t�m	��{��j�LP�,.Y�軝5�r�n)�����ݟ��Z�����C�7	�z�*Z� �r�t�SL/w�ߒ��C,���E4 n���
4�;�|_��C.�$���"9:\H���>A�b�H�^�4�b��+��$;��(��C��{��=�����i��Z8k�ŵ��p�bH�K�r)��>:�M����-��Ft�v�� D�2i�-�hK��ٷ͟lK=���-dJ��І)�ڞbQB$]l�������J����)�E}��r�1H�;��؅)x:���ړ�JйNh��f��M�I������8��Ɲ]nh�:ah�ȁ
�{���y �u�A�*4�P�&��`l��%tפ�o�Ec�1�W`ē�/]
���i��_��W���P��pF�e4<��i/�Q�y�����f�=���� '���\r-�jE�Կ�c���XV	�����E}6Q������B��(m��砟nΖ�K�Z
�bN�������l'|�u�z%�Q7yJ��WC�p��d� US�&��.�4���&_���	;���X�Ew;�R�2�$�Vc�����I@{$|p�V��71\��'%E(H�j`d%�QZ�8[��0&̹!2�������wU	��wfXd#	i��*)&���޽�&\u2��q�6�
�њ��r���f���4Sh�L��p89E�=b��� �d�R���^�mL�����d׆sq5�$�Bp>"�8���R0nK�S,@ gʠ���
#�Ί|ڙ
������n��R��b��))|��%�[��Ȯ1�B�����KM���~xp�
�#Ҏ~�abn2r�(�u��&�$fN�$�t�ĭ��W>ڃ���8�&Z� }i����.�t�����\Ud$���T5��Tj��5-����������jQ	�@�d�{!�=a�H�8$��J�)�!G�����*6P�DO�w^����{J�CDU2=6���o�x�Z"�nVt��tv�(���~�s]ZO?�\�]"�W5���H�������?v_��m2�8�x`5o���!�ԙ� ��?pN�q�sd<��p��k�'�]Bդfs�e:h��@B�B�EWǜ���y��u�!��.>��]��= �BT� �̜�i)��O��ӈ^eŒQ�ۅ�_(}������i�w;�����!g�V�/F��U�� Y䌃y�������t��S�X���(�卢v�m	��!�G*��!j��ǀ��Q�ʹ�p����4Ϝ(�S�_��vX͜ɬ�#�Y�7h���lHQ���ާue^]�Q���M�6{�_7�Ъ{�8_^��w�{昵���#��L#A���c"/�U!�F��:qMno;K��bSs�"�C��
�
�58#���D��t�{�U����1<g���������$t��0��4l��R���N3bg�t8\뱂�uT�1�e?f�LK3s����ZW�����-'�%��I�Y^rү@~���������s���itc�l��� \|Y}O��Fh�ֵ<��#{c",������A Ya!u9.1}a]~5db&�t� �p�NC�,nF%�(W������O��"�^0���lY�?��4�#Pʉ�L�#{��Oi�J%4�{K�9�����:�$�s'%�8��&��{V��Km?btꙆ]��U�C���*���q]Cج�W�)�Q��r�ٴߺ�z������U$/�ʟ�į�k Hs
%��Ev��V,8�u�5��>�YW����N�>֫��99:����9<�����1z��M�L�Ŗ��\��+�9���:�/�4��I3���E�ز�[���7�l��ۻ��P��}3%�����Q~�,�y��{��(��D������7�w�B����}2VqgG����H�K5P��Ka�|�w.�R]��?x��O�*r.<���6���ywݼ�FuD��'��}��懈�Q�V�^X��l�NΜȡ�bN*��3�I�M~�ͳ��]��&�I�z��4��1�;%v0Z�Mn��U�v��ow��ą�+�}:Ld�
l��Y����_|5�W�&�(�9���D���>��n��-�/��d���n"I�c��0B'�/�J#�b�
�g�3�X�pc��Z���s��g���@S�b�QIa����ĸS?a�.w���Z�kQ����x�w��:nCX��y-���~�/G&֥Ӏ^y�����▿92s�-҉�.u9����i��,���(U�iu`����B��c�4��f��f��0��>N�כs�I���gF�]�h�G�����A�m����X�Q��g81c�D*svR!C��Q���7�A/�rJ��1+�"��5��Q�PH�ͮ�:�19y���=�ܪ������[9��bjN�Rֱ,��ix���)+�ɒ��w'<|s�)�6��_�<��SJ�끓z������c�=e"ɥ ������~���|V���_��38ܛЄ���ZNhX0x[��Xw����@�����qD��y��2� �Z^@*�|�e��j�1��@V+P:]E��_\����^�Ph��AS�̡�cQp��������uF�ُ��9��94%ZZ�q���)u�(��Q�܊�@ H)*�"��7��r�W��;��^��M^�t�4����<ff������9��`�?���sd�y{u�\8T�s<�m5��C-�cS�-}���9���uw�M��u��4����P�u6)��O> ��C�J{����&���C�m�gauQ�%u�(roƤ����-�:�aZ]9Ǐ��u�#���c]�;���_{��SDBIl�N��>�����B��'?!�஦O"��fǇ���U�o��e@��SQMU�fc,�]Z�U$n�h^�/bم܁�)��=3e�q�hDՌH�Go	UZ&�p�ʉe�����A��{}iS��Kj��&t�].o�Q���;w�OhQ�}�@˴��e5"�J�徖����Š��^O�Ä%m���W0$+�3C������LOy�5�sʈh��$p��!�z�dŹe��*I�#l
���>��8Y(v8V�a�|��,�d�΍+����RD���� &��ң�z1d�i�+�rሶ�l��W�� x�N����Ul:ה)��v��^�'�v�G�L9�	��ׯ����^���VFl2$h��-�.�d����쁉Y��n������]�"��zV������=��v�>�����Ti��V.L�c��6�sb�3��L�\Wa�R_�/�z���ƚ_Hb?El�2BU�g�.����>8��.=|d�\3�;¡��ky����o���O��$�2O�W|������v�A-]�*.&�L�J�5�z�(��!��z��^�7qۑ�w=M��VW����_������`� D�J/�"����",,ǔ��Hz�h����W���\����(:����v��ԤB��I�����E�.���o�z�=����懲h^�?8N~5N׶��4�"��L�sq�e�<&������u!�󄏔��(k�X��4j�y�X1�Q��A�^.,hi1���NqS�s
��O�a���a��KVF8|�j����g�����������I��U����z��v�Kz.�Y0/�D�C���y�:�Z�,�p����7�B�m|�t�4�3�����ɜ)E�8Nݿ����_���v��K�vM֥x��/�[��Cz�NTVrp�g��������m�0�Jt��6}�.�+V����E�Y���o�1��k��]�޳�(#�H���[�0��D�Վ%M���+ h�*����;�(��
Xh���Sdpx2߾�i��̬\�	�{c6�Ԉ�G}�|�x(>��Q6ާ��z��I
�hy8�/O����X���G��7����ɩ�c���Fg��3a<�\���D*���F�-����Q�kK�x���\� �x C�kq��Tf?���zQ�-Zzl�DCdq�P��1�nj�2���f7��No;��so�3O�:��Щ��Xd+<L2�i2|Fͱnɬ�btH�>N�P�K��3}piK�4t%N�A��)<�S����I6m^�rGմ��'�r�{�Z���Q{Hܔ���(\��MxW��yuG��Ɗ��¹�nY~�mNui?��]7��ãO��?�w�n�o�Jyq�<�����㎼ ��sY�s��=h�$;��9蟁*V�UR]�Oړ���?��N�i�U��pXɐ��tkF�����؂��X-��80��'�̽�����������\b�J�J���7�:C����ØL���l�>a�YiCB2��Ƴ�����@
�� �zt��*�]�j~!��4��A�S2��,��k�����oAwd�^;���G`6�%9}�����mhf�HD]�.V(���៚���?ȶ9 vH���2E����% ���b��Pw��F�զ�\@�d��>{��}fVWD+	h���{�����q���u����[⨑*ѝ��^�b�l�,?����%��IE�l��D�I�B�fڋeK�?T$5��yU�R�����AG�CT�e��80p��s{{��k���=�˃M�n����W�0zJD�W��>% 
_��������4|�B���&.O[��+�{2�V>����i���bՀ9ޥ�?9�g�!I�G���2 G�:a*NNݥ�_h����"I���>�D�T�����^����@T�ň��B�+G�\B���f��)c�D/�l4+�(8����%��j�Qe�q�0��X�P�&�{b뗘J�O�-q���+.�M���S�\0�L}��֨@bc�D�VSA�{R~����΍��Ӄ�7�����[��:�f��b��UG�;t��v�/�uم4tP�h���_Yi(�ˊ�Ȝ����d(�������������G^NU���z��hl�w>_���d����ncf�!\,z�:��1`n�nB�1���T�f���5����� ��S�c���P�Y��K�8ߝj0��QwI�:��ݑ�����%2�p�<[n�eGNr��\DY/��H�L"ap����{UG�M��8g���J\o����?ȷ��h�I#,���UGY,G $}����_J��D-�����������œ�.�v��n[�Z�^,�<�����/
;1u͟�%�?=ȱ�+o���-Ȇ�d�w��{�Cτ��[h���v�/�2`���*������l�_������zx�fzDSSxcTT�a�%�����jm/�A�G2^��3�W;��=��Vl��$��hN̯R�~�5z��q��}�:)_��@�m�<�W�K�ɝu����HE���A��)�;�Y�����}�U��P�@�O|c������디Z��S�Ν�O���(�"�� �ǿ�3̪�@j�Ϳ�L���iR2���0ߊ"�U��ڟ�BS ���\ʢf�dsf<'IV��w�suF�����1<|�ں6�78�V�5H��=�s�cu�6�:��В����m[�.��r��c���?��!�=�w���	؀�2aZ��n��ވ�x:��Y��cM�9~[z�����O%n��&?����Ф6��a�E*��jN�h:d���"�9?/���yg]�2S���kzR8j��]�kI	DќB 6���T��U���Ā%K6͛�ik�T��a_����M;6y��Ue�6�$5_�PL3�	�g/�S(�L��/�Z�M}�/�����K	1,�59�B���<�(ߝ����/�B��|�sڰ�T������P�6�w�r�����{f�+�)���$��Ҩ��\��|j�_�3F�8�,��AJ̴��Ք6����Ag
H�/[+���GI�h��
��:	!�@�.�5qQ �%�	l�q���H��4̈ ��)���C��"@t_l �J�N�� qdk� IT�I�[����?�㨝f���}Zh���n4Z���b�V����$4�a_X�?bc�W=��	6 �2��f[>�K�n.x�Fg��$�Ow]�#JT���I�Y�����\I�4�y8I&$�K,	����Su��6��y&�^�h$��'�|�q~��V�ʶ@ )E��~E���(�]�'[�z���N0sſNhpBZ�e�s�g���e;���P��M� m��yߎ���3�B��~*=��B[=������`a�N;��M09-�0�i�O����i�S�{{��Y�f^P~��Yo�fkġ$-e���C�t���k!8�i:Q��`�A��%���W���C�bG�D�$%�:�R �^����O��;������E@�t�ۍ��p`�U4׷���q�ݿ`H�����$<|GH(?s����}���w�mf�4Q��F}jB`��]b0|3��;�C]��x�p�-( ,/�)����j�yY hHN��o��ғº�LF;�ś���aϜ��	L�	��tW=m(��`p�������Dg�4�3UJ(#k]�O�4��n�{�Yd.K(+��
�s2����G2M���ӳl+<�@�����u���o86��h�4d�l���=����⼶姒�@H[#Рp����2ū�*��X�y�&!C���>33R���*��R��rAV����:�=�Z�H��Ǘ��]*#Z�	��ş6���Xs���B�)�0���#�^o�ܔSq�vU��1Y�I�m�pJ��T�:i�qק�1���A<=�M�:�S�ɇ� ,�
}<�c<iĽ���P�'Z;� su�1Rx,��r"!�C�f�QJe$Ÿ6�U�����:�ݿӽs��ƘUk����6n&��|3AX�L�زn/R#���Q�\��MuN�6�-Ċ]yfKԗ�YX����u�?��ޖ��Q₯���7��,�2Rn��L%�����Scw��!+ú�{���;n%o��6Pa!\���5��� wF��@�d��O�v	7��C�j�ܶ��.~�k�gTrٓ��v�8X7��Yml�k����9���Y����������ϛ�P�f6�R�z�t��ō麮K4�������ʯ������[� �6IV:�q�S�$}�f��.�!HG��Z]�CO@�2&�ؕR8c���
vs���aZ\W���v�0J��
A�I��ē:,���W�z�o���&O���<�>�Dد�۲�Z�'�=��j�������U�25�^8�	J[��4�+\��"�[&v4HicF���7>���	T;�� ���:�o��1��G��ż�5c��D�����2I�a���M���{��le��Xs�ȃSm\Em'5���ֿ��^�$����\�޻2�yҟ�� >��7m��bR�S�)�����P[��F���#�ֺ��#_����S���*iK�[˂i�KR�ss��ƌ�p�k)Y�N��2g��U5���:�-����:��n�d��f���%�$t�s�Ԃ*˥@6����%����a�����O����/�aL�U�Y�5 �Z#����I.Vľ��"dPsZ�'�MǞ���;dL(��n�x���wd~'X�.�Օdj��u��$��D
,��o�C�/p�ѱ��L��u�i�~ňu6ό��LiY����dU6fS����&nC,��-t\���*�V(A���D\�}wI����]���l��(��y�y��})SB���+��A�����C1�AMT��=�V��eP��N!���Vn@�M���az`MK��c���8�cϑ�s��K�@�f��t����X��o���P���9��6��oF+�K9Y��[|Z\cd�{��3p��n,ro�+P|�l2���a�(v�K�*pH����'V2�Y����u�I�&,�v���Pl����Z#n����F��.��/������`��T�z2ҺŬ䟾!x{�����C|E�1ę�lXĎ0WP��q��60�1i�|l	@��GRe�	H����i̤���[����9�������+�Eơ �l���Z�7�`[�rW��[�ϪߌX@�G ڀ�V�TG��\�ۼ�"j��m��f)�Dd�k���b�+�6M�砌ØCQ	(m{�P�;��EqJl!��Q�:I�,��\u�Pj=@)T����\�`kSpR&CE��2�X9/s�Iq:�w*-� ��o���hk!5dPX���	��*v���L��!ٜ����C�M���b\>�=Yd�W�Zy���,B�Á:ލ�N��{�O�CaT��~y�>�	�:7��&\�Y�����d�� 3��	]/�;2��\�t_É� *2�~�������G�qȑ��
�J���;V� S��4:�������c�_36Nn�E	#-���MdUn砵4��Y��+���8���{��f O�J"속/ղR;.ʰ���u_e���j`wV��� z�uEqc���^��g�O56�s�W���(?_eIW�`6��(Rd4�l
�R��R��ɩn�b���(��b�q?q-M$�+�F�����¹�U4q��K���뜽���c&�Tbʷ.�G-�r~�w�Y��&F�=�8��-4��_cB"I�fn��'��rD��h�p)������h*ʜS�Z�]�8璔.2�0�.=yٟ_Ts(䋜y�0"�����.���Lv�F��>�7�W�?�'F��5O�1r�:�*��^�J߷YZ�S�"�x��4�!�eb5�m0�T6a���C0�(GZ!Rg�˻��dFW:���J�8�^�q-�I��H�}d�Sj��������J�[���`�n�䷗�֔�8�C�~�q0�����hcJ��;�=M�����j՘�儇�	�G���D�_)��(eB��+