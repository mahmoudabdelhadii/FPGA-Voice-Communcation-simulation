��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��,�y�}�ǰ�=4d�H���`I"��W�`r���T:tB�T4D�m�)�	1��I�t��
��8(�8t>s)ו�."[�漆���]�~�]��;�O(1#5�-� 偙O��QZ��~rL'�x[�i,mׇp���O�I43��4d�,�H�����SN��d���3���r��m���̨T�I;uj2Y� Er�*p�Q$Gm���p�V�`�2^���,hz�<p��l�Bxt�5��s��\yq���#�@W���f:m��T�	,*�񞭋����_��㧋l�	�\�:��uGd��PǷ��N�I��_����Tuv� ���us�(H�~�{2H�:Zor�Q	#%�3ˠ!��iS��95�,?�.���/�F�i{#���Tp5����Ҥ0{%���2vpn���X�����@l����3dc�ק�3	�Ed&3�ZN O���z��s�yxӡt��v*}ԫy nj#��lc��m戭k[��5)�A#�����8�!�]�Z�s�M���t��w�!��'ÒE�rv��Ϝ�c@<U��\tq+��&|�&X1)C�����r�A~��B�&�����s�:n{p��͠R�X⺂L^��R����c���f��J^?��ܣR�O 1�rV���:��T�4���AD����˩�F�w��)Dm�O�b,�a���1$��c��7t[i2>�ޔ0,S���󧇳Ϟ�ᒨ�-��}�!6��Jyv�醊�^_�(�H�(y^����o#����X��3-�k\8�M�T�"`R�DF6ȕ� �,5�;Ҭ C�k���1\������k�t־9�}���� ���QHF��"��t�9 ?��{E_�7��!����](�S��0�q��w�9��=�i]�1�GʦȪc�W�XC�|�$��}q�6����zf(����լml�dz������*�eLD�*�,�m�]ہ6����D�Gw� �g��' A��)�m���b��ӎ���o�6ūvO��=�W�������}��	����z
��z�&�P�K#�^Qץ�_������&�)�ٺ�u#uD�	' �/|�qf�M&P)�tL�x�?�u�����ҽ�����*c"q/�\��YDl2n֢�vtX��Q������ǰ�6K�gVL��ο��Q�������-�˚e��"gb�_� L01�D��ثU�8-��Nw�@�$[�>V,���6�����=����{>G6��v�����φ+Y��	�d�A��b<�)��Gp���k�(�vWu����!5Y�N�z<V��Ҩ�Z?����)�JL����q�]~���/�C]Sx|�b{q9^��ib�bl)�:��MW���SHC.+��G�~��m�5��%^&n/z���Ӈ��~m����O�Js����?P��"�� bfDF���;7~!��)HS �DB�t���;<��u��}sEԕ��)�!f;�f�(NB�>|�R�k^W��ds�@sh%�uY� k:�4ܣ�����d��d��:�$S;��P{�_��!��b�'&��A%<�ޝ�\��á�r�2z�iS
AM�����W*�}xH9=���"�fDm���c�y�����tW��hn3�1�T�e�R�|Tz	zPnDPW\�7�DɃ�K�ح��}*�ט}����d���&�:4� 'RH��O0P��<��Y7DiaRΖ��.�vI��p���u�|A�L���42�)G�ZT��HX���uU�F����Wu����_:ݪ��2�!y���`�`d�d-lE�Sn,�5�F�����,����Nc�U��%i?Oh�%#׌=��J��ן~���^,�X����iAAuA�q�@��^�:��F�,y�齸��Sz��X½��ל'��~�4jNT�Sn\��E�'v'�1o\�X�P��I���>p��lr)���0-���r�r��@gY�e�Ցx�����Ӯ�}�}.��o ���:Fi�'����ً�w�|��|�`ь�e��!���4!�����B3�y�F�fh���î���~�MV�ET��ɠ'!/L��Q�e�*R"ؒ��� h�n~�.
�2�շ������/7AM�݋�GM�A���f���,[o^��'�8��9G�J�O�Z:I���@hH������q����5y3��J�M�����Y �`�9d�,���s����hAƗq�ht�	Q_���L��Y��-ѕ���jե��r�׉�;��D�˝�Z�vm�W��a�6���3K��lv&��V��6!��2����?�����A��}@-�⒫]$f��3@�s.q�'i���▣o��7̪����0��`[!z4ْQ�j⥀��BD1�{���V��g�؂J��<��,���<`t|i����D�X��Q A�ޤ��{^(Tv�y�3�pܶ�_@0�׿O��P���
�'��&3Q˙91��̴b8��O߂��f?���Ú�ly��V݄K� ٪J��r*�vr,}l��24�ňYB���yoFY�%yϭɡڪ��U�Q-����C���I�/��b@�1Rڧ�>�F_)���C�j����_\t$���9��1���m��G��584q~����-%�8��E��Vt�\�,cuȳm#�8t�:uk�����yPQ(�>e�P���d���t��hؿ�ΈfMH^v^�Y�+�]��h/����%�]C�q���>#߳��v�DV��#��Z��w!�vq�N^8�9}7�#R� t����.��}�5�h�w��s?��Fܓ���������j��y�6��	���������G ���+�p�:v9&���`��>7��C7w�$A�M�I���.��~�
��	ʂq����jM�?��?���R���7C�"�VV�zC�ib$�jڰ�V���*��3;?��хb�>3�}ܳ�\Q�DH��5��5ZBok�!|nΚ �hM& ��:�U�Z�aKlؚ��,K@�f?�;,����L��O֬,�\�1d�nQ6I�ּ*H�T�pb�y��6�?wOA�J������ӄ��TA�	�@SC$��
��nLY&4-#�l����Fl�������18�����s�ɱ1����'��֌��d�w0�=���C<GѰ�)@�>���N��Ӎ�Nj_����
P�
������������?\#g-D��Ő�p�1]\�変.d(O�O
�B2:H/�9�k�-�g0��h��
G����.j����y���^6��
Ȭ���_N�HۙFƲ���jhn#jA�ÓQ@��)N�^RI��3�墄x��B��¯�� jj�\�mz�l�)ӯ��{���RӐ�H>�*��x��w:���/J6J�<�5Lsa*�f��� �)$8��eI�����5�+Il��c�:��B� ���E�@�`ޗ�g�Ѭ��њE��L�NH@�b�"�r�R��>��@/��K�YJvn�h<Q�<�h!����ߟY}��ajvÏ��/R�0s�bF��Fl4!���$�l<V�\avR�k�8+��xk3!�t�I�ۺ,�%´3m�Tq ��q.#X�0u�AZ����i�6����ra���HVq�c*ZT�
~���^>�A�˙������&`������剓:�9�*��|`ѯRCU硅���C��m�c�w����#��JVv�G���.X3�,�x5׻���u�5|I��Q�:��]x:3X����f )D�Z���:A������3l���a���\�,�{j��ǌஐ,�S��W&�ܑ0ҥ���!�,��p����v�{U'�[u�C5�n	]?�����NC��=�����1��K�w���`��2� #R���.�h0'R�}4|�[*�^���d�NAj�}��9�l�w/����"`���q�dF���'� ��` ����"��&�Y���A�P��`=J`�`va�R,��g�-�E��X�nkȜ�
�-�`O�*�E� B#4�u��b�!�e8�����w8$LaE� x䏬�Kݡ���
��[�p�����i��>,��SԿ�C:3��_e���w���_9X t{����nqu���ա?�\�a.ث����vܷ��D��1c����~�P!�S�H�BvZb�?�����;�+�!����l�a��3�Ҡ,��)	
�n�)�Y\]�E'fiѹ5Ϣ��T`�����M#�b�i�Q,���3wQz�N�'�y�*�;���s�] n��6~�M!�hf@����^YS���4{���)IlkxЫ���'q�˝�p����\jx�Dm�o��/p�M���^�&3A�}��7w�C��vE��8U�(����q
�(-ʍEy��s�q�!��F&��C���⋺���>����#�K��n �T����{4ޖ�N̅H����-/�/v��+����0��XC]K�q������"C���9�0���b_�9.��c���Ӗ�)�WN;!c�ٌ4��b\";)M�5]���ؔV�e��Utա���1�u��
8�[�Pr�Ě_�Wt�����4����^�(:�c�
':.-Ʃ�� �N����b��UA��_5HJa��#��fߍ�E?S%b�����cd������Ufn�����'��cpbr	PC8zMLe�l��r\����ɏ ���p����}As(��KN�/��R����D�}�NG�1*1�{��m�v�T����Q�B����~^�����TBl��'r���~ce��~M�(�C��\D#[*�g��!*FT`0&��٬��P��?e�#����׻�?��5��Ẕn#��z�?sa�L
'�!P�e��o�q�/�c�E�^q;kl�0�]��Q���v/_�8�.|���B�%�E�ZnrD���%2Xp��ֱ��x��Q�h�s�����9q��
0#��691b�p[ ͐EAޭ�G\����|/_�L�:�/��n'[br��V% �>91�U�}���"8��`�Z
���F�ќ�l&�i=�`��r"�M�����%;��&����$���:�.���`�h�Mű�lL�>%�F���!)Up�������	Y��T�1���=۔j9�����i���(3)?��f��%�m�0}�.����.��uR"~=�Vu�ΧІES�	޷�j���%�T�>�H�F�f�m�� �0x���6��9��o�N�T��1��NH<����������p���p�����
ƹ�A�5;i����6u�Q��ws`$ζ�:v	��l~��X:�vFw�s q�cq.V�����([��B��9�&��]y(v��J��y����Vd��| �&%�L�Y��Ef����QA�\�>���A�?:�-_�u���nD��l�z�B ����������D�Wh��)n�	 ���:A7(Y�[�B���Y��}ܬ���o�	�`|�$х�W�_����JRW?��l�(�aa�Y���=�ѳ p�?��M>G۹�D풂R�svX2��JӤH&N�+-����K1]�I�K��g��\wN�쎳4��½.3��W�>��\��9~}'+�j��R����>`�c�����Şܽ�.쯗�ϊ����؝	�: 
����!���4L�:���]FE?	�`g����8Ҋ�'D�=aC��r�(?�
�m�>�;)�d�&[�-Ly/s�h���p�b�y�]Cc�6M�ml����?�.d���yv���\��<a����JN�U�Č��ȳH�w��欈��^�I�;�����O6������?���ֺNo��ù��lLw��)��R��D+y �tvt�ez��yقV(��)�ߨ��=�ų	Z'e:�b�?bnE�1��&�J�N���Ќ��3y2�w�Թ��L�Z��0j�8~ُ���(>N�BN!Ί�D˓��rƷ���������-t��YV��)C|ڗ?|E���f
���>�� =;0��\��'G���	�XV\:�g�pu̮�џ��#���f��f�]�1we���e��� ��d�a�\��#�P�Y�������<c>Hn;C�\fI?j[���6YW����ف�����v�i�|��*�%�n�v�46��.8��Lgi���ꗻf��	I��/�[C�2~��4��^5�l]�i�pe�W�����fѶ�r���ɖ�`Y�2�����v8NX�tI������F�-E��v;� ���*7$� Qp�h1p{ylԒ|\�!��/�g �l</ś�F8&��=���ܲb�'�j؋n��(�Zd9}���%t�3�ɅW�����!�3"]���+k���M?a�l�ջCEy�I�[ ��fq���$!��(�/��	�ė/�z���*Js(%�=��B����a3�>1K�x��9Ph��p����d��<>��M��Í�?H^鴱���1�x?�S<;��)v��|QqqZ�ƃf��=D����e�f��n�M-}'�3���-)�d��?��Q�~dH� ��1���t�iiZbw��j�
%s�V��u��Ik5��Ǖt���sȟI���.%x#~�Y a�'��#�!Ǵ�C����s�a��[֩��͚�]w*}�>�����/C��@�CBI�d:V��t׮k:9l9�D,�bR��/Sy��2���-j�I�.��
���E-$m�/���S%�*xU���3���Y����=)��Zu�Rф�`3��.�A:��M23�`6�-۟�\W�ŀ�r�?���$�4B�;�&��M�A+�Y���Z�������V@>X�`X����F�:ڙ=iP�퍄ђ�M����-ӽ�J���L��e)�r��os�|��p��_"�s���* ��%��گ	u�8h��R�����a��u��1���Z�9�����j����=.v�V�y���AI�Z�%��3Ol[�2�J��`pa�e=�7� VFK=
��4���7iH���K<�V�Z5V`+�k^���'(gh��s�R�*n�t��7�ߜ���
�$��rO�s_�3�h�s/�{�T�v�L�N፱�@Ìp����w����x3��H� ��]��\󪐧r?�2��!S	$SE���=�3Č�RF�צw%β�_�v�W}~ԓ�#%k}�h��HP8>^�'�gW���Oƚ@~Lx����k�@ �I����ό��u����1�{\A��c)��r�s젣6�lp��$dEp�+�j�6K��5I��\uO�f�}��g��Eh��"I.`�RZ�h9'>�o�����)��3����^�p���N261�
�*�x�7���=�ra��!�c��Ϩ�f��E��	�j�#g�|��{�J���h�m/<�إ�z���y��9�CO�Z��R'jk"�{�A��O�c#��F�P_Hg ��z����:4$&Q�A�.�N'�E�qo\Y�=ؼ�q���N�YH���t�d���kL����\���D��C$��<z#�^q�b9ĸ�`zN�I<8�.�Y��[(��<��WA?Q0���ܰ�Z�3��԰U���.^-����;�ѯ4H�9����B������i)>��\(q}��q^IpZE�����P	y���3�`��Ae��z�ҭ�a�@���w�C��ӳa��,��� j���~%��8�F=!L�\m���<���&TꜾ��lޣ��߄<Z��I��9=��"���͢����Ox�x���i�԰����?�����%�'� �PV�=�������������O��ɚc��� ��5k�F�
������o��"���� ۊ� ��ޔ�,[�&�\M�D�����Ê�U�~�+~8��9�ۣd^P�0q3�ǖ=]��@�׊�!���Ř�TJb��R�X���n!?%��ݬ^H�7A�"��E{;�jV�C�����ڥM��ä�o�8��ϙgӎQ�%G��������5+1~4�g�x�Z[쾙��1��q4O��3o�J�^t��T끤�l�Z)�3d�.�W���Q���6)Q;�5V��W#/]�N�ӎgl����ׯ[i��>�	�&�E�r D�D�Nћ^��9������@��]\�뽪L�%���?����/12Ŭ��xʔ��yɖF�̾��L�m�C�矦�.�A �2>6�� >��z��%n=�b\ATb�)��[���=]ͻ(��ݮ���o�W(�!n�(���` r�]�B�dT��s#��*�fTp��!$>�Vë����*��d��mW\\4��Z�&����NX�-��螂j:��Gv�c������S�;Z{�l��M�S�c�/R(���c]�1!�"���1�vk!�l���۸�z�B��a߄�:˴�`8&���{S�NFaA�h���Ԧ�޵�0�}�"�`���o��آ ��_��+:�XFo/0��*2�x�!gtXl�#	���0�ǭ���9	��)�]TW�JI2���u9
�G��ub-k�r,ɹ����4u��k��[ش
�!o&n)>SⳭtф\��^�.w"��oIh���ѵ�Zk��5Pw�-rZШ���ۄ����]��~��Q�f�S� �\�eMM
o�Dՠ*�`�
�Y�^��8��d��3��Mԁ_qԍa�8�|��P�c<k��A����D����_��֙z����[m%�ӑY�_2e0�]R���Y�g͕���e�ĸ"�B=�xC��,��d@�m�9�$���b����p�s��zuvH�z({*.Priz�?T�աR��P��l������NjaP�Z�@��5�
�����kҨ9>/%S���������~��zYF�B���L�K�~��&�?t�b���ֵ�Y��q��G�&sWu)P��;��{�x�5hEK��^����mJ<w0���M���4%�L����Ͱ�`�OC�÷�?[|��J�I:�zeʆw0��"n:r�?�O���Rt���]��gm�������ؗ%�}WP�T��P[�6�xS����λte}
S܌
��5IkS�2���-�w� j�Kټ�s6T����C��c��
�r(%t����
`J�R�A����K�z��@M����W��ɻo�(`pG�P;Bpk? ؤV*r7�ÿ�E^��r(ZL~R������-Q+oj�4�p]���E�NMq�J	(=א<���!���7��)�~Њ-�<��������3UqZ�1��[����&�A���y������w�K�{�WzmD�^����{�|!':_M;�NZ��c�)�谶~�Q��2���䅁�H	@��Z-E9G9�P�IT�mNuQ���7E��5)X�0.Ы�)��͓b���t�5���L��	�j1Lq�WgҬ��u�@�߻m��}�.�.m�� �)�pF��ѧ�,g�r���-i��o�hQ��a�c
x��\�;��T͂5��R�3�X�,��4<ϔ�x���C	頶({=ǧ�cy��齀��o�cí��o�?w}Qzg��e�Z{oR�'�Huk$�|����4e��c��hұ���bT��1Y�����5{�[�r�T�L�)n�á�R-�U�f���7��I�jC� ]����,���SͅL�zഃ	�1'�W�0W�"d�9�Z_�T����s�k%�s0�8~�]i�JM��<��VV���i��p�h�4^�E�b�y�4���)�$���`��c?`�朱�/'�഑x)�1�r�[�u@'�.:føj��Q�鬗-� ǃv{��.�#i{i�h{^U�0G�@�0�zx�����[��n���>ɇnQ�E�jJE`7/��xc'%�2����sF��Ce�#��q�}L�j)c�/�(�m�qf·9��GR+L��PI6p�׹	��ær��Ț\jȢ=����}�u��$�?,��wf��e���]u7�� ����u�sɚ��fO�,"���3J�<?���XA����1"ɋ!O��l4w'-�zfy;Q3dL>�5�%��$Ɂ؞�F�J�e�\Pd�Q��͘�+ԕ�"�
�c����p�_�'d'hj����IP��u�3��J�������J���}(�:r䮮"�5DT~��2����/ ����'Ճ�� 	��J��@���48BN�>ÙߛIi=?�:��p���U�R�?Ԃ��D��{^�>���2�Q��
�i�KaM�(���۠=Ҭ;�?�A�Y<X�"�T�Q��*�`����ҳ�=Um�L�O6X�h��|
�e"��,D�k�<����g_��mLm���f�xm�r�9r���\/iiP xJN��<V�^�A�5\!a���P=Ae ��^�⃪y�dM�H
6��g�W�ʠZ!0�9�lѱ��j�I7�H��� 0�;uW�1�M4�Ĺ�]�B�xq�@��U�C$�0���.��Uٙ�x���wP��dk5��T���:q��S�]�25��Ɓ�b<�����̲��HԿDUg-oC��J~RT����^����#[��:
�XqhjD���f�=uE�0�d��w�TT����V��Ff�wm�,��9Bp��-X��C�v��2F��B"�S�2L$�\K|5��t�L>�*P���}���t�7I�c�?�3�#���t=�)mm  ������G	V�n��ҮLU��mc�9B󺆮�F�������յ9@p��,]N�Eh�$���pkd���0#�lJ�PS�ș1	�KVE���xH�����_� [X���U�����j#�T���&��"��=��
І'�
��Z�$��]�Vď�"x�}�V�i�(c�j�H���,���O��k��L`���\�-��f�Ã���/tmUe��oR@Û.S}�U0C�z�ɖ6�T�qu��翽o��'}<��Qoȥv�3�˸���j.^X�'��{���^�Ф������d����d����,6�^1s�4�w >򞷊z���PN�G�[�A�{5j|�èF��g�����[�.�2�*�A!j�H�Y��:��'��j������{W.d% ky�aB+/��[U&�P��Mlh]I�+���k��֦�tNJ��/`������z=*T�8=�I�敇�T1!Eq$�+m�L�~��']r��E��G� ~\X�-G�A���n{��z�5�~J)"��*_�:��	�ѯ�����}�F���EX���J��H,!>�:�7��6*�^��5kw���p6_$��oG�8�4-��I�g��y>壝η�)�����O�_�z>x��_�z��ç�@��I�p����w(U��/�3q�=߱@q�^�
x��4P��h3�]�M���3�=1����s)P���d}w77��;��̩q�� )#̼�;|�a�!�$���y[L�������n�F�?����o�Kka��k��|H�{'�[Ǹ�) c�q�:��}o����!����?}����αgN�FvmF���&�)��7P���H ��Q+��:�=.��,}�ů�9�nF
Lh-1���F	�B�#���U�_҄s� ���/2��DU8��y���f_����<���H_{\
%q�\��Xc�����Tr:oiXNj���t;��j\5\,\��fPf�gn���c7Kڼ|J�	�o�B}�׵#�g���E{gu\����\,�.Rx�[�G���� �7���-x�A7D��34�؛;���Oq�I��V�f��&��:�(��Uǆ��vȖ��%��@�_�<�@���z^�N6"K�T�iT�H�O��(��Vb��p�v�UT�����wB�UV�d�a�l���C4�,����y���lXcA�Ukv��8P�(e��D�͓��o�I%τ��2/|�ʘ����B���!A8�4�R���G���m��V)G ��XӦ�v�r�z�p2*Asr;�
��A掊����7&��#��ٞ����p�:��^藀۔fGǋe�e�V�������:MO��JJ��y���V�@I1I��ɚY�Y������"Þn��1{��B�0�$n�l��'`���	F[nJ_��p��ry7aD��U�g�%��GM�J�u�T��4&��g��PJO�'��Y	+�>>M� �;�pfa��׀
�RG���%d#��U#zy�=�ߠ^f4x�-U�ٔh�~l2/E���)�_���9�,MP)$Q�C����+2�Y�d�sݦ�H�ʢ�o�.�:(0K�z��6U�r�<0sn��C�VW�;�w������4���tE�2D�V�E���$�f���	�!s��e0:i����9|�	q���?��@�AL֍�#�ɿ�ԻJ���2�8������L� ��Ś�t<�Jqʮ�͟T�Jr��
:UJ��Ep-�"�/ֱV���9�O�
�FHF�(q���ۅV<S�3�Y\p��!iJ�MdCPp����S(�U�%<i�2����>�������b&�p�\�Y��!��ʼکg�r�m�*gV�s#�>��j�&���t�fz�\%5�N�7s�.�v��˾�L�[�(7Ď������f���x�qt���l�ʌi!�B�9a�I}��%���Y�?}*��� ]���E BŇo�|Q3E2rHkw%��	i����1/�T���W	��D����=QA����$(���8cB��nl�90���4?�1�i]�FY
)��UX|`JӋ�^��� `�^fy��$�Ӑ�F��vK��胫�M��d��W[��9S�%��M�@��s��'e�J��P����g4!'��>����	V���K{��IJ�}��HL�:��Z B뛲̌eP��}�ӻ$V��������z���wr���z�Lm�������[��:�85mZ���qxR��V, ���)4��!�|�2��/)�.6y�=h�UL�sЌg�,?E+4��Z��6�y�XsV�wA�mjF�x|�pH��4-�jnK��A�d�(��蚤�PgQ�+!"�s�L��"+����W�a���-�z�B��(��h�w�����$Y�p�Z��_�d�)�S�@f����&��C�� ^��@�8�̊�7��=�֢���N��'M�3-~&���Q+f3׷�����QX�l_��((Q�Ӵ�S�ī���y�TW\����:@�b�9�m�K5g�Hh6��$�����<���#@Ԕ��1�����1}z0*	�C����2�U�_��[J!�ʿf��^���^x�H��/l|��n�s(~5h���=�BK�m[GѢq�|72)^K���~�:��Q��f,-)&��k�����Eu㠞�j�|��F�Fz%�$��ߎ�y��j�a� �F�ƒ[�̬V+p:M�@���|�_1S�슽��_�	n��L��m��vTgd�O7C�2u�?�Q�$��xZ�2t� ��=��+����mf�f��-��'Oa�ub<�^�rb��>q�W�	��;�r$ھ�5^�{�c��O��M3@�^�Ap����v˝`��U�H3�W��sդzw��ʿ��I�γ�O���+ܺ5Ò'�F�F�ߠ[4���A�l�D��dRV��{�C2i��	�!y\]�*�;�R#F��a�q����E�Ce��A���HQ�����h���/�`�R���s2"}�C�"�"�g���:��O:��#v�a��& ��,'��S띇d��{u���f� ޢtqd�gH����v���u{���$TH�f�toz̋�ڻ%�(Lc6wcz#M�]��iڃ/&b�;�p ��Hn�1E��v~�5�!����q$�I�`��e�]���7�F,Ko����5"/o��O�>*����kZL�
��I���T��e&�D���Ӕ�����f-����L��l��U;&2F�F�@.� v�N�Ţr��no�"e�ZF���!@/Yp��:�y[��d)~uT#*�v�j�.��Z���!,�!��ƾ�ɤ1UBZ+S��	�
H�o�GrM�&��Z�l����/?��|�ڐP�=��\��2�).mv�5H��z��c\��Dw�<���U�@���$(3ð�/3U�JXL9�U�P�`I|��q��)�۷l}x�����4N,�D�W���Z�
BH��/_V��4��_��m�����;���;��DRie��XSD����K� f\�����u��u:N�OѰ���Nc���w�L�FN��]ܸ��*reo���qĴ�䘢����i�`���f�6�΅t���:���t�MX𠇛F���@;��V��e_$�P���9�Ug-�\���Q������)�t{I'<��e�:V���+�L�=+X�fL��M8���`�H�We�3����0���]�������:�������OR�3]V&h��ǈ��ǲn(|���r��1DQt�36'�di#�mqj!�� ��^�1f$�F>�Շ ���Ղ�I�L�?6�-�"�GcN�n��$;�4�혤��xW-��t]����U�J�7r/����ϴM>M�͖~~"�D���x�AрZ�
X""=���I���8Tk�3��`�2�_R���9y64���y�cz�:�Lp�1�2�4Y��6���B�e�b���ǈo�m!"!cU�}���m`
�:�I���� �~���'���V�����Hl���=q���a���.�A{�ɒ�����.f�(��=��Y�<�|?�����,b�:�e�h�QG����D�6ѳUR:b�D�f�f�]��vj?���҂v�4�Pj{�֮%�96��{1�C�e��i�qB�D�e��?��v�t' "|�����awlV�.�U�B�u<t��\V�z�`	*&I�ľy�����'C��}v藤SP��޴*u�$`�B��$�C%�E Q��PUj/��dA�n�(-샛�̅�l��(��� �!�n�bG"WPS�>��4bT�=-L�ϲK�5a�:��.�¸>w�Ta���c�H�[�-w��nձ<1w�;]a���1�I�K�}�'L����w���9���:gSm��+��jzn��Zٯ�;6�z��p�ϝmί+�?d�le���Cu�ًr Ws��5z�
���X�8��x8͢;�"3���)`�e?���/y��
b��a3���w��a	���V�cL����� _pR����}�,�1�"�]��40Ԥ?B���}�p����!h�Q���ʟ�ˈ�)��)���%�dds`�{=6kDY�č�m@���t���r̓D��R����U�� �f���cy5�����h\�)���<���np_C�b�j#�(Ԓ��u2�)�G8�݇-�ϱOW�l�BJ:"�|w��D�YW�b/��}b��"�16��5��RƩG�h�4�=��A�D6�O��4g��5H����Ї@��Q��ӂ�w-�9<:B,���!� &s�%L�)�������)����.`�ohW2�|K2!W��Vې��4 q[wh��{ �-'��D���$:�`+����%��Y���h�t�f;[��5i�h�-��c��o���B�אַ�<�N6�.XG�Fl�k�H��ȂA���C�ȴw�l8)�#��k1�RJ���� d��v��&u_�lI�_�0�4!pH�Ax�-���/�y��)������2h�K$��S�g+1��5G?%��>ku>l���p����S