-- (C) 2001-2016 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
MNv4WzeunQ3IZWk+GXdWEhyiLuKsrRCLOmRAG6HfsbHib/5tbhDwK1TRRoE+LwE44Tqe7QNML0+J
7oHLvd+7+5cLjChU4ZJilHjX+Zb7Cq2w+ya4ikkaFZrknKftt3FeTqerHoOs/0IsYPHHjuGb88IZ
CJAMyyBx61fE5xDPtm12Svb8xuzcnQQgNNqOUcPy7IMnBdij1juRgWyWwT6ohNP5dN0BAGZAt9rQ
bno5aUfqOgW/U7L3c5GyvuMTdCjSCFom+uyFZ2E8ajlsaK+wI7yWaEsAGeXP3KJMQXqM9JoHNKIj
311GDrii4SEEF3TqElS1iK26kb6KJwu9Dtx7og==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 11328)
`protect data_block
hme6eyuC2P/wGK6qiuQoRiEQKfg1BAjY8nOfyHx3Qwlxakm/0vf0DAorscTGhwG8UCGwXG30SDW7
6t4eH9VAwJTqh2O3l0OYcIVAHJB5V7/SWsf/VTKmEJI1p6Sg/gYZDEDo9XIyf+TOAJOTlo97TLNt
Pj7r1hPAbwO7Ef2rxu1Rw1hqBSHrSqvXc5mj8AFECo//YpwMtwJAw6zm2CaLRQSpRcfUMqrBnHLa
J3V3hyBRSyWSrBqIdtyqcKkBJWUVxsSotK+gcw9oJEGzdmVnO2CCaMtZmbaAXO0GmDi0K03+4oXe
4UdsBSIIxZ/gl6k+YAvhmPwUzv1IR80Uv6Wz2sp0jw4+mqK1p67X3dsvRdmGwjNxnCY3Yk+FIh8j
5z3LnpCsdoUoKbh8NvGvXgi9Z0cTWa5elJCu3lDsfroutdrWaYuvAeyyZJkDonvx0+bhD3gjAPeZ
xYl0HoRBWKjeCkr+gkLlSxqEohiA8eAv3kJwSAaMaVseOwoAtkELrsNPRFVTLkmQa4kA4CTD5TF+
6W4VJyAonnS2sBAyPmyavoDh/FX/FBZCrOFFL5qtL1BvVlre0boYEAvanUnJELTkMUb+hvvgHhGm
JVYOmbPMyZykGT1JTw1afiDhkSHGbJgLMa4LW9kPrr/4rPMEzkL38K9Sg2VYBOCsWPhZFPSbCS80
oEodWeT0gc6xxkEO7FjAsZmrwItIu7rdpiA3bvxBAUmt4YLU6F0c8KZyHvtIfoKYAZfUMWn23sGE
5UrHOrUJNNVoBQLrc57F3kuncwdQh1kTZNjwGgmMlNmFVklGSlfxl6wXKWTpO1UpCZf6saOqP9we
EfMFol8B8eulk0OGKyhQCRiimD0f3+BxClh7P7i+jhZyY3MvqFEYwPzimForqj62qsEWEDl+cJyu
jYlctvXskooyFneEtSum/lDCdGJi/gSRq3AhZlSsnJOiGqeP8eFpyyQ7T3nEw52vmIMiwQtqIDYy
3XkYWjY5JcS1jR5HmXiz3B2ClkUZ3lHdO9g3w66yij5EslZUU+V1xV2yo+5DOWPRGXRjMzi64fDQ
g3M9eINZxsgYUhiM2/Gfjm4GyrWgpctrFBu4eU+TD0OyJ0RQhKThjKMJA+4bo0myWxc+oI8T/sky
RYVkCZA9mg9kdtr4CNjdTyEvoyNStA34sVQReL8ED48mJruN5bX4fItaBwJUir2qa3pIqEO31MlD
sEl2Fui9tIu9YvpcWQt3elTh9OZOxEKNM0qFuzFkz/bSyZhXWt73zPYwxJjBqG1w8FphkamcQykN
feK/NxxKBRL4f5vh9PSua9ada0kFgd83KLiY5BlP9mm5jZF3CSF/Ml2YQcNuBIYa79m7UhCaiIY1
lZ+jbdLFJDya8xnpkFSGHkHHu7ZxzJaDXuGpKIjtI33zKxlCEWy+g2WvhdSyci5kS+K506gWIobc
tNLEvD6cGelbBRiMqQwo04tRfsJwkYyNNOYBYIh0gPLVW69jjBnmxXcYPGVRVmayH7Bv6hQeaTeb
8XYGZlzsK8LTLSt5AwnvlCFw8wjhq/v5oPfAsW/1yTO5/VsdZn8KbjVYwphxJ39czSYJWj17umzY
wAbRHW63clXpY6YLnXPcTY9byubqcF8APB/Yq8gsed82nHTL4AZfkgelkVYRD6fjbLaUWaZg6hDw
0w+MRJJrNnP5soELc8GMqWsPPWBwMGCMR5+x4sRRDEZmTAMpA/75YZ7xnze9r/aSHpBnIC8l4fwM
V8sSft5D+j8y5oLk+zbc7YcVWq8vq0Cxe296IdQGEElKAF1/VpsS4+DXl5WlaxIv5T+rgE3UiPM4
joCVZmA2x4kxzg7kqVZyKhy5TipyAS0RFGdUICsiFMBwzDe2W7RR/mjMTuFMc+EEpNOwFeX11AhO
LMFoPcYeyNqDensGSZGe4dsoe5H027BFeOk0IwVR0X2gs+2bN6A4oew7P2qSZ7sXYxk6GEe9omTI
kcH47ui87mslxSmQN4a6VztP5GmjHzTIxzXqJHnUF9bttsOtF2z3n9GFPCfR+w7OulpwUM6nycFi
pQJxs0YVGXSWDbBqo0rTBrD16x4tDLyBOTc+4FfMyZbzrhl1dViDR6XBYQmNPTsYr8G/PKPOwsfv
y47jdVMRHcynUPFTTFWyfI8eR0l2KREUgZj5VF1FZSDzFuPdpo+Gl/v0IYx+oEvDmFSfgWGoq0F4
jydxd46ZwX+6LkdBn6eHvg1H1h7ggR3rR1vdqn06uZIwfURpLfr+NBO5JRECqmFuCdxJ/n4IAAes
wyQY2pw3zD6oeSxM0tHtqNXnGcTQZDZNEMPzDk8JO1hQ9DHrMIaVNsiJcbx/EWrgJkUoXvSUKQI9
z30TjQuQBdxwoz66zdBg7+ZkxbBX0D21sorpYp2bVU37ESeo7a+coH6UsN8R5H0cWH9C5eh5wzy6
IzwDyOo/eME/xViCZaXJQ4f75XKLjmQQSCnM8HKBhxmD/YFo2Ut0Y/VbNAIuoQ9aekNcBjNiS0r4
jUOBGQgNyzlGI//RXNf5+Ua5FZH4Tddc5HVQwW7G5DKO17UcZABr8tDusEB478odf/Pls26eiIu+
OpfSP656XNwbhaQUTrBQEf5OBDTgBvebZxRWlz6U/fTaj2/pWKncmEkMWQU9nvxg501l+G4dMPyn
dnXYQ96CBb/WH+aXMY4fiuEmDgVCVWjxOFb2iUzGGZ4dgt8sVHBe1SljFh9S0BUdrAU7TyXmGfik
665sjZKRikTM/PkS6KXOOua1QT1WwCVRjMZqVZjVskn0dJQr5KVLLE8BXK7DhUkIDu4Gjy1zfXDh
S87ENIqOSEqTKANqia4WM9vF8tavzoO5oNHKxb+HyYaWlab56Lv0vGsMVLEW3BKZh7Qrth/8hYIY
rN1nuuGtPP2yQ3+ECNZ1QSHER+YmELZa5v6PZ53cHkaeuuuB3FWPQ2HfwV4zVEY5xwZTiVHqyop+
XiA/turu2k+NyCB6dIygU1E8ehjxyaQGJlYqJrQiuzWRvI4fuvAZyKSrW0KiGpBBEuNudAn/6J6I
S/eGN20GqAkj1I20QFPUNOzYErzG7wHhq8EWX7yyWpbcut0hyyC35sXHwm1c1VZfcXpSVHDqEcND
2c/s3EPzuopN2b2E7IwywX6nOkMdNAxRowdgEdiWsLtqS3pfmjpejWUQPnqoAlaszwJ2tmbJsc7C
p6ic22IigGy3JppIBamIMzDktihT863/6Wci8+BD9v2hSoUX4WphN8mFx7LDmhjBtza6zyIU4eJ2
/DRK+Q51KEb1omiTPLKBtXQaMRfC9D2OVWbLA8J7wF9k5oS07W7WbFAJQEelp23XWFq60hEtPXpt
OXMey2uQuOPIUxaHQgQc0sA6G9vTRGHp1hqrknZW2246j8wpJdFV9fXPuIYZZQo6Asp9sFxcL1cK
/sIuAyIkwt1YbOaUiEJYJ0xX+jDPCTd9isQ2BiG5+YoL9DT2eAperysc6okjlZLv6YhE5nscxNp6
MOayhLq9B63cKRUaxfOPnO9KKL5piCb1/zv1fYFqYLc+DRAcBAZnq/MwOph5GHH4h1yOfuqU7tjG
HWGgMe8uEJacG8pY/MNPABO64kEaLMYSnGAz0c5GOZ01gb4XQH+ztUL7xcRd7MY26kDh5WkT73Qp
2TGolyB514+6xd+cvIPyzMMjJiwSOwc3tTO6Q+TBjN/cTyOP7nqcwf+m3iJ3IkLhPpDPzspcuask
lORTF4HJMUjHbEj49Fk02Mq9HnMCkMHbZTZfZh/KPAqvl2xIhS74y9ff3spMIJCEr3ipUH+2sh3c
OEVJtE8LEj2XHHJIDKGEp7FY2qN8mxnsRrGOE9wbWXdBa1OTVYHn/kW0k6Co1aEbDkY5aBZdixDX
F5gwIkjwx7L84SSZiEAmFGYNIShghxbsYZmihHNglt9rQJRhoQoJJ8ZgGfqtlpIdQyHbisr0Wm6A
5U0+yrJH7/UcRn0UdvjvJMeVGVyE8etuDQGtIWHGCOEEJtEW86OvXl9I46oqnqkPLu1dpxQjcXuh
E5Keicnm5gXOdp+tqoYUk8ieRvaX1VGqyA+lQ+VlBT6yGJPQVwGCTgtvxWPGrAu9Mgx1COsDn0MV
EdZINmCachVlefTc1aEsc2jlR/eQxyr+5LYCk9Ecgji7T+2uekMsfpluI4JYtYZ/Sie6ERe+6g5E
SUjeN5X6nU2Ihuqv8MctkWP0droawNhHZGtnMJFmDBws9+YwJTaf/5nazCfJ8PSv9X9vsdK0kBQX
sqeG7RKfo6GS8D9Y4rcI6ek1cd5GqW6G5mYUJrxX0ZHBle8VFjBmFTVxUdokmwXHuPM/XyY8wXWi
/U+CXo4321mH/eAqLWNrWDkjyELI48DF7uZ+ee+nIIPwCoa1Twp0wpyuGZ3H7vMKncsumgVXW5s+
2Ah6N//EP4eMJbB90WhrHP2BbQpNHQwatLwkhKFvkUjzNS5HJYyBqOdbfxMH6cTKccNHjIGetbwF
Swhj1+dsNeKJztBlh7PF4jov6wFG5QAjoZs8khUh1mNh49YShL3xxItJrws3dD6hZvffMLOWboyL
Z6h5oSMtjnkfvyMO535jjZqdqhqQX7BTWDsHQc3SAMC6aQEKKQpIjKIvHwpXHFMqjVstk7lR7Fwi
XC8j2x/AmO9fWK+qthoijquWBj0iTzj8U6G/Pq7ecxPMzT4qHrArAmpDIIcY3/nmYMcn4X7QU+mH
JI4Amqn8Ti9+kExDkcunFVqPpgAlnJIat3IuoqamYEUWEqJIqhnr1yn2LGoeDyKeIzFvUDNTvvC5
rq3atRpnlJQ/ZXH7ueRmY2DE1JcolPvEc6UswBeDOHyHROd3epoIwFvur9lzeoAxbg0bJYkaXxNJ
TDM1nNrMMmO/1Gd1gVjxBCmp6mjGjmNrzTeyC2s2NsIchO6OU/w25IdfF24va6TjZqriHAEYXF++
xaZUXmfE6glJx/rMoYQvjxr1Ec1O74QWqfiEZkFAklFHV6iWzz8yU8091NA6QSK1rWEFQZkuI9F2
Oe1Pbm6EINlv997mFM3HGtbTAZ38woMYQzyTH9niy+XwCn7o32HvK7aUjfcIY7ALdpyXqqi+XWys
K7q6XTAbaosDDfTkEoKn2cbJGssefChmtjmuIctpOxMZA97YBIGUTwIcKF/Qj//PxYntzFebZYpr
KhQnuqP3D8JNoZGsBEbNlAWxXUJpLOCzvY6TNqiqHH46OplJmF4DLeqBz64wB8EscxnYEiN7JzK1
NC9yInAbTp2FjsyHKzsE5fJalp1PT7/+Mpd4WbOjdz4dlS08zS1eDf8SkjMoaHFX+HALY/qLdu9Z
QFgt3IxI5P3brFA5J4eS08+pgHAU34m669UYKpIZiRAAgpAOxMFVfVBXRVwnbBH4X8Kuzw+67sSf
LgZzI1B/3wtW1sylMKxSrAExe0QMD8452kraWUCW9wPLTcAqXuHQfj9FqabBgQQE2vrzcmlC1qjT
YNmqKutpKTgBZNti7/0gG06FpGnEuwTlnyHj6qNpvivcrSsxt4lPP+FcAhcyrdWGbIIZHsNFd4TM
Sf/ozwWMtmjwFTFZdPuZIPKV4NSUyLJmbW2I/DfsEbC8hClaxnAmOpiGxr1j58i0VoHP03OZz5cE
cS8j60bE1yIWSigOQDq8LwQ4ptzxwqG1PPz8WZy3TzFeKYqdgTMkP1egFq5b0Y0ClDpW/I8dlnV9
kBw6yFv8FoSpRbe9l0zGZ70RNEJsCRAkKAMFUDr+yknp5bpbVIpVk3DoChfa6CGfba92R9jpVE9G
ktHbQlEub/6L4ePtUNFVD+sP1NopAPyVfAFy7c5shYkJ5GKydWUPBr9qXBCnIW4UovRNLH8ye5rU
Agc2wBJeJhyUZEOOvH/t8IQdoCyis7jtqJXgL2q0NL+xMRftJNveXCTN22Rv3skTEjyklIVocUkD
7Okf6g0ArXO+/isAfDMJOJbVISG32brT7gaz1VWLim0znIHzQLer6a57K5h0a47JGrximpmJy4G4
ToMFMdJZg0In7vRopZOSniwc/zx/JFRSo0SZ2AGZXL8RjKLEC5Y5R2ASgaixrnSdEZ4h8SvdVjDH
98Yd03n9KQCn5cRiBVGJHZ1lyEJ+amLKj9aHHa97s3ESdNAy+Pv1kO6UWFTrTLVrawvCbMFnaSjJ
Gq7srvXKsNaWZAzWK5aoNH+032QDl/U5xS5uznj2cX45DQPy+0tk9Q5o2JOJJCRIWdvp0lNfIJFn
ya72jlTdqMzXfK6nJhsiGkAxcKz6wGViZqD7pUjoHmSdAKKOzzimG89YTktItIQwWAJHdu2hNiZw
RkxdoHxbC43PZwqebmElODBCzA7LYEsmA1uMN1+O5HDl6cdL4hHYC72LT5zpqIxpFKAriRP86Q9o
m+R2YG8tsMckQpw+rWa12eFXJhvmhASFgcf3m7xd8dLa4PhOR4LBA3K1YigJ22htyZXkyr7IzGik
aZGuTnlHNEbbtqpSl9lhfCcVCJQXsJpSzglDAd5OE78j/F2rEjcFqJiSmIw+xcaxus8Fu2QGA7vk
VPungkWUrEb9lKFONkcY6J2sXkzrRH6/r8sqe6dOHArIyQTBI4MwpGeqJ4JenGctLKMq+sZBlk+O
jgwosOyk4b+IJexM+A8EYIMQp8eqEyGMW22yoJ18g08jgjrGZBXsGZaIu9zh14Pzttihp5RZ4m9g
XfAWcZQ8lM1sY5VRL9DeTrXVXvPxAyx3Cr7DeqssUSR5G/0rXslrzLDOGes1JQVoTYrlAlN1jnYN
P1PaVr2NKNtanc52wAWVMhEXz8P+ovKUYaRxtBUqEe/+aImMvhUBME2QBaxZDZN8z4gS0UGiiSMW
qbLFxuap2ulSx8Ga5iJsX8gNnAmVHBXsixlJdSlrBX0/vNMzsSC4YTS4saltSm+nK+yZ9ztwK6VS
iZ11+l62x/WqCIQ2Jct8w5lVI3i/upG0PyBzgGcXHTIMLcaqpAPaqh3kJTl6iln5BrCwAtrrrBAY
FHby/tf7ry2c41WUaAi4JShC80ewFY5/9dI5ztAD+sL+Pr8WL4gK2FcL+dVLzYkguwhinwh5lRsO
WHWUQOo3XCxg8YB1++8KVWn5D2oGSTMNcrFxB+Igf8l2IXFWa6vx2qcDWpMewDJF0HwjtVByozs8
31F5LiHvMyiHk3YivFGDQ6iZe2HTVY434rdZDVp2Z2/3GvuPXMoz43IrJsqxYS4pPPqAi3iX8umT
Gr95uEhfhvl0rUCNsWck8JR+X/mIuz/gImNRO2esHzCHqVXPUL5Y2n3znst9aLkQJaAgWDXyyX0r
2Fz2Bm0pAymWVdUv4gysc99y2xBFNCdyJKAjGbm4jVZM+u2W7HF26Vmfj0Bu0RvFGE3pxrq+Jdoe
X0lqita5WZt/XgwhNEz1HouItMJ8kcE0a2tzxFo7cX0eeCW8zkhIMhlhA0WnRoJc9aNeuo8fCq1X
mUoXsjylAqIV/X01nwYOew8L32lzrGQpTTcks6i6L5MIg8Ks2Tq94/KwUaf96QIRwpBwm70Lxr2u
y9woykdHiTRgLKeSRdwOepqO2CLBJXFJCtyCpNkJgwAiOxkAsfkjJ6KVpekuVIr6RnDH1VN/VaxX
cj6kxQjNitKfRYNOPWuj4xMSgZ4CNpgkHR3OnISBRKvfXmVnywW18URs27OSrlDot0FwD/DGRtTl
PgrY1x6IAKF0CuRTZt2fSw61AyLlHu3CvG4pVcEOH+ONw1qaYfOUf1aGlgH6th27EQIp69g1eBcp
ufkW6CQl9cNyy5rEkpi5qHBBgBVLzphMOihH6Jruz2Hr2Tx7SNni77yntW5bYCQHFdcUvR2GFATL
QLa0rZnCHw7oaw0BtZqrMyT4gfVt/eJxnLsJ96VowjZsv3HkRuOTXHXsM1Ri2b5vEppTQ0Gur35o
QXFnBbal+5n8+DpIfTvCLQx0tyK2NO/IzgyCvdyZmgRIWbciWyPm4IoQVH2OQX1tepQKLVoJXryq
KD9VB8rWqawKCP+O1VG14NQKHTBN8sv78JkOj97FqKIpaBa+PWFMVOSo6kV+jSjAkvwri05o4MmN
Cc0dJAaZieftkqOtZ9jDFUzIqnztaIqphlyMnLk5CFZ753m9Bnl2r5e3CG1EUYXAPDYes/sOc9iE
ZatV2Xn9ZYtFdQNksQ03bscd1/NMLlS9d8qYnoSnYU4RYhR/v9bzwT6u9+eYV6HzT5/CjWbS2cSY
WrvHa+CDHx2B7a2gxF+3sjOl5/O98AqeoOExRaFBVAzdl9CyWfYk0Zz0u2WO+qsSlLTZJfdcY5ng
6JrGL0HBg/WAhp1rW6DsFJVhZcwS8uuRLSKHO7IkxOXHvym/bVSfxg3Bff+yliP5sSC4K7ACuJpM
FlIcJaAHv9jJDIOUHIRcbpir0KHRyEbFIkcMQ4vTM7O3WGkuKV3NetMXjtw2gFKywL+d6aBA+Ivu
d5doyht3PiMnJ/T4q3PBGQ2ejlzyBUYV1MTrJ37npZ49Qb4pj2FSCUy1HZiBWRUzHfkozZXuy7Fi
1jGFOE7yow4T8eVBBcmkFuVwR5iWlLOKomVYfqGe4MEgfiSjh4u9txbv7Y5JNcsKiWPHcadPLtZy
zlel5ZV4ZbYwqP6xG6l8n45c98wu4YwqxNmnkKJe0QkpgqVKjtQEiX3tm8b1oJ9Q+TqPjOmyJAeG
k/ZarCg5auBJ4qUREVMUJLzTesIjHA6SOVzVqJo95TC6Yf+AxHE6YwtPMKUetbtkOxj0PhVsO35k
x8zgLO0qwHdGuXSlLG1pdk8L/oKfU8vE99sR9JBrWrNzzd6LzNWHJsHG01LnZ2Bw6YWYB1x43ap8
pp8cTbt9nD9sMMpzVB2DhdhmDBM3uMUfC9mEZphRPIDQQ2jA+OlAb/L1BJqvb564xAbe80Db5vdn
mLkQKPQFpeimUpUuK/cFpw9rXL5naSRo63AzDquZFVx/+D/kMefoiF2wtVDJfUKb+UayFOri4r2C
evdTEwQAAYG2J7VDV85lFXWkfAh4QG0R4nBEVw7OjzYtoSKPxq9HHmK5tixT6ZyB2pgT3wq1A/Kx
85VCr9G8y2WEpc9SJUYEvX2PWoIL7lit7Zr/Le+hZzHUdG4ORRLAGjUeqBO1XEQA8aUzQq3Xd84/
Xjr/zs4QwGtEdvpEc+ksxd/FE2hYFVj8fLIV7hldqUdCztbFpEYcu3R8RlMi7BMGglomfu2C2U/d
wvVxDd1vhPBjfMc4Kizc+4J18ABAwXwc6B5thmIqcBy9my1S6GC7AJ37Yvcj1VfQM67MuRbEyvdu
WJzz495P5QiHDLDxbrznIqwA2LWyVePNXLFLipUCi77HwvDeubI25ce2oEmf00eN2cJskE9M5TRR
rpLT1gXwEFylVL2BAIaAdtwP6XuJwCqrbpcA/KH6yE4yOlaro0Mj9Z9eEJoexDlSYj6pCPfKsDN2
tzQZhZ6W90nq9yvNmVRUXxHz2csZfTBcuLUwv9u2kktdNNfMpuDDjkEGAxQ1S53GvUvYFJ94f2+6
Y7OKULoPlyI484GcRhMKwdZECUzTasiFvQNP4+tXn5nQ1aY9oANowyu5X/oDw/esIWXLPFdLUIbx
wOloRuNAMr687DxWS9Vnb0//gSQdZ2+T8BvCF9PUC4KVfGpy8WsfMixCxRXHiVGWrML0bAODqDsy
LHAXGAZd87G4wZ3sAjUBVevSTsypqy6Bvs4Hj4ozpG2ffQ7IEmUmNf9z0o5Nz5Far1dIBFMZjRFU
RLidPWONHlfcN6dZLTa98s7T5oqeil5XEzLT6CRlQwNiBiYEgeV6OTVmUgvIzFDgbpdBXdslPQIh
0fJcTwXiJaelxCtP06N7RjNlsrgR0iRZxRs0DIWIk/l5Tc8hIOeDiqoaDnaw51IagJcLXA/yee/e
eUBdBaC5qwTooIicAkRnW55xB7voaAh8LN+E8quGfyRrDY9X2T7NGOafJHcrvrLHIjuUGaTNAxo8
xi/yD7ryiYxhG8g9lij3y2YwkfDrIIQU8iIRKtdh5uIdGcmwzABovEaUflB4fVFGwc4PnFLAQ9xn
8bcCfRrxDpUAY35kHXmijpPBj9FTPmAvqBhLFtV+JrgKJt+44xRxtz2iZjDPoJIE3bCbmfmNjB88
i2MZRVFtgwuwOSFH56RNU+bFssguqgXR1fIzPP9FK/dGLFdG+sNOGegRFZzgEXprOm39Bu0+TOIF
wKW3ibrKC3xab+Dp7/53bVAjypKREwcHnBgxPI4h1jVHP5og7NcMSt04NcqhkjiEdxQ0DmDiImv3
gZjxLHaW8Ckpo+z9zbpjFbgEE5n+jfOYA6tcaJ3gcEkWUR4sBzVoTdHpjZK0oecNb2P95UDexE/d
lxvDhNU+Bi/Zq4ezMkjHyXpLnasuyYcXZozFuEdyGux9nTS9TbV140vgUZKrHIuZ2kda2fiINhKi
vXpINnLoPMXEawnBdlNjBtZVGFES0vMHCaqZGWZNN5nwO1SzZsUmibgm36nBIgV2X/oCReL5pT7r
GfiLWams7PPOaYK/wYMKo1hzRyLVX75XI0In4kSlPSAF6nrqrMwdWolRvPEGfXMo3ecfGkIJc96U
WTeGr+67bkiJPeu4/1M3K9fJmvRiF0RLJnqFHUWYt9veEXUfdrGKHO+YjpdJX5ymvXVsA6RMVGrO
uH9qQkmn/P0WV+DoyH0jNjljVMjHF6duP9+5NQ+OHsOx/1dA2J5T919u5vA6FQderxk6zAATUrP1
fqBV+Eht1uvviocIjLqaUA+BYYNJGd/yjdueG+s4PDEeo+EcFFdf4ShdMkGxQvXVAr0N73eggZZ2
blMKwWwKCOwrhb1uGrqeAvSEf0TZoZ0IWHPRWMEQn5tIAk2ozq+3J7oPl3LM9yAHY1iUajDYC5Qj
9uM6L26S8fuGV0FpbYfBiX9y3d9wzacxoq/eKHGk4JqOqBDQPhTy2JU1atV/y9eETTfAyIif1IVd
HQ5+BayCWpHQHAu25hVTDhsFF0wqNLR71MujzXOgJS7JTdig2UArL9kxqNZ6oFxmmobCixnqobhb
xqH1FWW2fhwFeuHw0ctP/ds6SBvwO7EJ/5JrJfBcbC/OjDthW7Y4AEW0wTtvAf20R2EEE8wodigY
RzR6M6KCv88NsklywacDuHGgv8N2NX5jKqmY4b9nIwTo2js1XEz8CTShC4ialWjeu79oCMrzk9Se
PHx8kgsSY3/k0kU6XgODsIbirPWYZ2m/Z0ouowpUP93qGu8AoyEIYDSuqrn9vWQwEUVSaXwngtgm
NsHQh06a4GKhLoJSqhPFouHd5YMlBUaXlSjkank8u2JMHd8YP2oPnpM4C1OSVa7ChJn6uYhQLmOI
jnjoVDzj8waJrUTuESUt2F9Wdr+3BuwHCXoVixAOsPJtsd+PN0rFJbOQLWvJ8DuNc3kD13otZegt
Ddqgn1lqUrE9uiIZWN91INwN5GcoOjRolQHVpDwkFTgyjS3DzR1mj5fBgND6oS30jUz3/XT1dU2e
1T1wjTjMB0wQKdxOiRdYtRCLTs97CSc3UZj0oWxJohHiozuOT37flWirriQppvB+hSYJCflPtThB
4clbHdf3qBQ2qCDbM5Zwdnmodm75LyK9UkVcdyDA5LAd2MKr4qsFovshqsXoBt+WT03BDX3oS+fE
5LKfQuE8KqJb3PqXIkYDoHD6yzzVZ9biub4fLDWuXupbvLWtR2WH+chd55qZ5JDQvjXXFMFvga0B
mIFrx4r28M0IdvHhw5a1nIjByQJu5Wlnr2/cLhVkmkZL8yWRUKmdIUmmhZ5Q7gR0nVHwXkY8s1fB
8U9oHaytXhtJxO8oOcO6s8szC+bTdzeUXPa8MDIWejnz0rrAoiaYocpXw7eiSHlnHK5VHff/ME5a
b61p+abbgTfbx8RbtRTKUYIk+iJowQvlr/SN1GXt116mnY9vHoKu2+n9np2h+RP5bkfgKqPRt/2R
JTdyAGKZHyIzjLo7/ucVfzWwXscMETUI7KzkwcUfO/eQnV8ouCA+w+NEnSerDc2FAs6v2MZb9I/K
E8ZBXwfahakOEKAaVyXBcQ7dpn+2pVnnCzmkjSZBjVFXGRQ5HuL3FmPG9AGP4q6nlYVdR9MicUMN
2bBwp6RPbrBg4et6qqmPDIng/dIx2UKg6Oi4UpZnkfOF23XI2c+2/BSMR1BTUG1ghwFEsB44BEYo
WqkKQMMLDgERYA4Yl1JAdHwbu2mt/2xzfpTSrsXa0PzzecBnrySY2KmJYoCHw0nN7MtlARTcUiub
Xaumknu99HsaUIZz5FAgA1Ickx00ocVCLbYfjOBT5eyfQxZCaZ2dRlBBVu0geCGjdI+JCFsD5S/F
MSnvutDvQOQMrhtn+R3ljRDDh8z1BvvrH3Ffwxo1YedYl758IoSMwSQYxnItYDcfbtJmqdYlHrIb
Tp838br+xI3Ei47uQ6X2QpnkLc67X1JefyIm5GVtmm9Mhl2JW8ZtbTODjYjh31jnLefFPRwEYSnr
0iO5Lewcz/4F84HULmBuMD1WSTMLbgtU/04wmVrMOo5Lg5Wg6BXeibu1blnr8uzj+eZ81yHC3Nio
K5AJOXvRSZ1AcxtNxAFaCCXrJOSJGMTKH0QMG16QWTghJYMS0G3hMR4BEYvQtrdf1gg6Dptbua0m
5bK4ufOxlKVLmZ0boIV4tBGjkHMEnFD7tiW7yOyrSgSVTvPwRIfeCmxOane72JFFsAxscDx/YmDx
iEqo3W0fHobuMt/y3K5vBLTBtGZbR4A4uc/QHMo/GlFYOYp2Vf0RpxjDjD2esQB9deAnC01Ow221
vh4al0F2T0+LlELaNqEmgnZYk57EoUiGQ+ESsG+s5ijl377klvKyUgs/8SH26I0sqVZ5HrR3TiMC
37Z1n3kXTNkgHlZuB/o1zVGBsG4jdCBFkZMsSd+yR7X2o7tVn8CDrPCxFKhxzzCyzidhyTjMskC9
zl+JfP7pamOblUe0OtIzfUeWYO5UCfGaRCWdbdvKrbEYWIJXEB9Qw9Q6Sgcb1AwQCIhyuhqmEhi3
j8YkMb5642TZQg54SUSkl6J3RzUc+XCYdKP7o15Yqa/z3RCNmbfkl+H/jzb8Alum+1pGh7UrK0ok
i4zKJOdu42k24KacyPV1sVZCcdIKc7psdr/un1SBdSxP+m1UCrc+OSmJAeFqv6O1RcTrKnNk75pn
zpriEDlBI3XQP9T9L/knahXFdMGPw1POEKvxlVDNPUzMrtaLepX5W8NUgmoQaLlYXwKIEmJzNV0f
bo/gJG/3KX4/CPaOOlfTU1GGrOkQjmoOjZNyzjJ4Y3C4PkwYrDt5ncPsxMDbX3ctR5WQIOZCvGdJ
XVcCVIPdND5rAxUaOIxXaOJ49r6f9R8mH5Z3hxZBFAiu5fLkPwH2UyNd7gA/aC9BRI3hD/UpJJDB
49Yc/eZciJupTqFKlrevokNC3AbAa2Wx5Cwbjsx1If/hDmQNAp96QALuxW4LoEfIu4440THlpRI6
Y5li2m64TgPs6mNFCPewvRWC9TQTDcC4tA+FK1ic/EGP4DGtB+Iw/NSqQlITqeSDTSXdeIsHm8x3
xo89XQUi7joKXINfB24r/wWS9a+3QdZuSzSc7IWB/od0Z/dGi0croZqkmFAXk9j7zbLWiKvNDIWV
PXRPHu5nXqqzsvUTYQIPGrjiuX0iH7Qdt8cRNNs8S5gKB57M290RZXRq6k+sdYiKJMlAeEPriL3x
2RZ6WxrFEaTP+q+Wn8mbGPoRyggLF4CIRtGYgIvzNE7eQWkxb6bH4nVxZLGJPTYRfxI4mAuW2xTT
T4vsd59DTM2dMaVdkcabnGMsNNA8hFT56kWSI60kcX3ZV8VrU9ra3a5WxblYaQ8352Z8f7zyX5bQ
QdvuJ/2BDo2XMAr3vOxEFLh3ZQddAOY/Ta6jhTTUWo2qM8aULl80K+FzvjsGGM4N0vAjpw2L8P4Z
vu5bdOOzpcWejXW6vUoNLvVZZ0nJYDsFe2FWWak+L+YLyZs8H+PaeHAPwHjLLWDUV5eEACkqcHMB
tvjQYAmASL0clQcixAh1mY6S5Cmqh5sZMXGCm1Xvtr7TEQ8tHxYPdCIMKF4c6k06Y0cyMVCUlGrp
JqkDgRu5c5Xyuf9prpBJa6QFg39kH1EF95MbJSlOfXnNIUWrRfQUFVEmFLO0xzo7zur45JLa0yQH
PlZnvNoVqzDqmw3PfypRnmIeVPW484tpeGMphllW0ysFeVeMC2sBuezwf94L4K2H43kj+TuYmgHO
WO3T9aBgCGEVSNhAv7+sH0y03k2eQFji0kvRvH+rj0S7rzihfow5V5ltK5c8gY/85jONJMasi4SG
q53EpG/sQsAY6Lj5SQYLW4znJCwt8J0GQOKsHiU0LmYE8fAgZOs1b1JXrZsJpyuWakcGO9E+Fqo4
awHvIg8EJK5dDJSqe8s1q+gQbgRP7ir6wT1KTw7w+ohGi/bQ17/FquRBEe119GAfYVCI4Wp1Cvlm
yY1CJtozHAi0UZ3NrX/Hvpud9/t6S3KBtFdMFhN9qRbdS5CCEJ1VlZFOOTVndi00VIjDEq8GJtvX
nusc59QDrzeGfGujxT9x1FmW9ZYrGXfIRllsjSQV3y4pDGef8cliLUz7wsR+aKpfJ00p9ryajI6l
6BFXIi2qXH+2SVpH5oe7e/8SQPkUs1uYErdkhBtS9liLNRzxRE5wYVb+tyewKtB2G3mmXCidyZMV
nOhNspcxsVbBV+q6aMVmWDC1X+iz6PhQPVk4V65f+Yoal9VZNFjBSf43e+bCOtqUvRymwHt7biPi
mw5IGjko8Sfgc2GMXKAFpViUyV98I3R80HDuQiWOsyMlBhH5igyE1yjjxF6H5EncMl7RkLrhQBAH
oZSPYXyIyOSDKrC3n5HD22d6/v/CLKs/tCpNU0iBY7I6lCv5PTMyOjNG8yQNyHQJ8+x4KMAQrgOB
LtEBLb9Wr8bHvgug5CeuNnQlqQKsv0f3/681F4d+pL6ePFHuJjWkO341x1Nld5OBgjJ2LNtD3ICA
opWhQwsZAJ1+k84Kp1ig27plL6Yoy4Xd4GC4CrVyAktRVnmirufG7KciX+lLU/FS096Hgtb/Ms0O
zV+Yr5LO+/le4QLRC57Eo8odamprUU9Ld0N+/ichECSzK0pVS8/QQt34
`protect end_protected
