-- (C) 2001-2016 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
AT1CRr+boQ3qLWLvk5tSp6Npij2rOOQDirlQluNzjX4ItL4+dHfGWkqR2zAUos4WbwskO/7nPYI5
OziaONCmYqldZetp0V/+ORMDm3HMpNIYp2mjRIg17KJ3OqvzASEa3iM1BltR/QBQ9rwNqs104/eJ
A4Xqv1wZmScnH2LQAwdK7WWNSZL/QZPyWclE6Cg1aAnk5+s0AzF2oAPm6I35+uviSVPphsywt2Su
Gv0CfykIWk/l1c0WyvZDEf7oYVizLVA/9WXe2smq5Mp0kbblgXo0nqGZfm8o8iahLZQcb1UZT2xQ
SiQFy3jQjoeaT2h86wpdxBcfmVfw3vJmgpbKfw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 16224)
`protect data_block
pvIDNuO3dGMEnX+8hpBWjjdsLG9kn2UCwnf01JPWMwDcDrZZRibHU0nejqXh3nDa2uuL5sHFO9gf
H+BLb3XqU7tdMLhCuW3U9wdWEou6e+xv9r4ll3G1FZKawyBNBCpjCrJibjkjTQT3pDwKuyvufiFk
Oujft3QAMNqjZbdrQpCvHMfITRjy9WLRFsNWMLV2zsujlBY/9rxZqT/GKXcOg8nXqG8RY72BjUO2
vwuXxxmJ2Nz1z9ANeJAm4DsqVGOicwD+Z8SUhjAAXcKI46i2jRXBZ80Nz3W0F4U+VoHz5457jbMI
rH7Tdem3qze0KOdsjotql76XwJLs9uk120W+/B5/SHR24bZNERpDsK/MjdT/NzL3yRWDjUA8kiNX
9OlGU5dVsTgH1c0G1snGXXe8XtFx8vFxQe5R6EaYI9HJpwYJvXRgjXlZup4Yg9SDANSsvOGu7WC9
GkzqrblGKSOiDJaWtLdmlt8HMBVtDhZzZZTozRIZ4VTksuZS6syuXVySRRLX9vbsn+ak/fx6V0zS
urrnrKNyQmVl1YQGOIuzftRKE6Qf2Za/pQRlKtgPbEMUk+8Pcl9nAQGb5gGHUbV77KhmgufIsOsK
4cUrOdzIG9shnf3YQWlhHoNgJx6Ak7immRBfCSZpwvdnFPywINZsErXN24Tzam8MnS23T1O4Fj2W
ECVN2rKiyck/yO6gyoKBrxuHDxJfpkiyjac2cCL77f//zygHvlMBfpfZ1B0ao3+u8vLFhqeYgWrx
wOdvaMUeWuh+UP0nmewfFxbyi6f+f7E2R9yx7GoyOYdNPHkj8UGE4HRc1QCKtvFp2YxVJq17Vjr7
5101MnaM6VdYye38zQTVQNgCagFeH56tp1tqOJ9qBk/WZXYjKZTGzLehNEexcqEp57hbdjK/nBEA
yG2QhwBWi9fWtYSTsbjcSJprb2EOLWcb2fyJ0WDMtZn9V/cpZdldmo7WFFuKAGG04nfWJ8TmmiS3
CbN3hOMINT0X+QMG5XTRcFwN0a3Qd6sredYTPcwkhYadTKnxC4R92ywAClOYR+WtkqhIYzYR0K57
I/QsudIaB9b2Cur2rCQ+bu4fm3l13QAFxoAtdKTUTwt2ayPz2vWVKQL1wMNRM8dSCi7DPFMEvJJ0
YxT6YzAQhPvXn/zAkqFY3OMZyjQja5qI/2sibhZdI4prA5JE0UxQIDCHOMYxa1bZOvwYPJ/pK2qc
nRH1TlxP5PNrsCI00RobAfnWT6kIKQcQsMrTLBnTH3VxL82Y58Dq1e1iuMXGXLT9kZI1TjbKrHV9
daBLi+O7f4ODwQOwLVRX6VbpmeAjC70RrpE4LrAig5yxTtAoFWSdEGwSKcue6zmzuaYdjZ7p7Y0J
8snlwv6olwFbOCPmGi86y9XsysrvvYAJRpdWERLRStuhFx+XjfQR7xdBKVncoZlCcwCDPMr5t158
acZZpYKgDSRYwIF9LcIJl5+mCYRSUWexg/EXyAzrQnal0Km+dbRYmnCH8oA7sAuuCyq6kg4+2GCE
53jrXv7JbMrpZm/QPOquIpUjIGVw2XEZbV0MF4o9uoPlchr61zhvuyOpiI3VqWpOdILtAZH1FxMk
ros6VEYgpdYkBbriULbI7sKSCuWs4FD0WYmdOVE8P20VL/hQzW0icQtCKjZ3UzQd8zvdrRoiMBfD
ZRY2tHoy2G+4MWQYpGWGK377Vei/Zp2SvwVovUhhGokprHlCMYihFcztey2gNbbkd8CCJ5Ksje5K
2d0TXuIrvQerefdLtRwKZhdC/nHHf3yH0j/RxiIaJbgZ3Xjme+aNkajpp1CiCydNL8+ECmtz+tg6
rtdYweWjwsuKXaoawzR3mt1sGYzXfdf48Y+CVfHXM78yAT2ipeGsmj367nHCcU3U1lR5ydc4/llz
VzmVuKpO9kaak5VxxaITO30hE9BXdnziSbKCFNTHKOZI+SMdUcmcVXvsHwDJUCa0IANnDd4xis/k
G1crby9DEGCxAvHK+Yn/bg3U/kki3L4HnuLtyqgbQobl6ox8FuQQDiIXICAASQ9kgUWP98Q572qn
24j0TZQAzUYda44zYLLOT0B1QCV1AR4F8GV9vJDa6f3sMhHFG+9r8g6xEVd/hhmdCjEYsCzI4ima
+Yu8akBoW5XSmNM7J9Nu3fkNhdUpQzaeJMoMFghgE80fFQkoI8/jVsZ2dxEEpF1cE+dntDDUqRzi
J3wlPzbvQVA6PFjtNvQh2ZAd1CKf/4Qpj5nq1311xA1FY74qBl75FePc9AEOYsCxG5peoukK/ZQ7
nsx5Si5YdGCz8wWSk0z3MeIEJGJPaviV5WyQgQglwfujFWTwyKqqvN+xxiaOsA4pjEvSKPXA2QfX
UidBqmFF4gQT/mxyo5tkcFW87RwL40BVzgwxlTZCAkr7joLmU6NxJnTkgUEfunHk7wTo1kMG9R0o
3q30AI3IET7eC6NfA4O9NHWlvBz8IADs/t46VfCt2OxevoIvFEvqmzk9gS0F+TgTSi3Fitzqev1W
jZL2sjUSu9U82U/bERt+MOMfO55eKbwcOJRgeyzkRuZPVa5EgzYl5m3nrEG36eXdohTC93/UzPaQ
neeKUT7nrRb16flVvvfSZ0xMZrwC1eGhbh/Z/Tr+y/+Z5igcDE41k+/ERGuP8bStqe7UetaMrIw1
afsl1wiPyrAsP+/E04QGzqrfS7WhIXEB6vgBzeuYZQr06KY6HXUSm9m6siiTIpZJxXRFeawmaFaJ
skTqxvATmqohZmHDOH+hzDVZJjbLkTCPl23B+GTOXCvXsOJrcyyduG4esVYyRVEVEIIZjl5kPb30
qkvVWHIbQ2iJmZBBcYpeqNvoawXznjqe9oMb2ZXByl6zoRKwonAteWuYoUF2tKdTI8wqzWyWasyD
785QFIX0Qix7912FjTITh02x+WjWlI9SGYtX/JUh7VClRb8ITECMmheJrDDL5VjMgXxMYadKmAPk
GXyjt3gE491f0INu3YP5BB+9cL55zTiF0aLI4nT/1li9gL0vjUyBXlaonqOW9TJIt3Vb9Nk+Zpq3
Eo0A2dOmz1bP6u03DpAb0NtDpbHZswMuXat40wvhSPx4FFgGhO25UuuLWcWug969th8+AjNEJkDq
ESgW3fCfsNTZsW409iORNHcBUpZOEfCPwE7dxFotCpgqagPZ27U7BQ80cWKuUhkjzERd3Sxw/bof
7okJxnjkLDQcNHg+OK3LrPO/VCj/LKk7r6NksgJJ+vRXcLTfzrPPe5BsuzM3yTeDkTF3/UTp93Ho
Im0DpCC2rIkN8wh2NlrM+XhCfOGJDUtWAfer7GSLvTsWl0atsT2V7MmOG1DYVREEMd7zD1nwwfIF
wxnQ89aBSRLZfIftviPnb3A8iwhIb+pwEPBdZkJXZd+WyDnciQzkgtp6SQ3U2Mr99CWO3kIE5uRc
5ZKlixGUVPCCooDbkzUV0HMvCLAz8cALN2a535T6VokzNtrvLotlCixFszngaGy8C7Lduc244+Es
t2+OnyEHXK+TwjmvZJLbK5QZg+6wAE0tRtSADr+Xm1zZegNTNZkFKhCoUgvDe4l79MqinAMmPkgX
OPpXt02tkZUBxmNieb3oqwgGi7CFYxiM+Pg93t0/7nLj/Zbwczm/9FnjkgLCviZZUayEDIHtcdeG
nycTtii9akp+brd2x10hdGhwoMWvGb6junbcTPXCUGyx5KrMmjMQL8FVK65aZOaW501fuNRJFJkV
n23b6HKMpNKgVmF/upqpiaTLSZ3Hch0ABFJu3y9Ah22rD84cvhu3bdQHjBQDB2Oha8xxHNRVkENu
JWqMoR+seF8CunycXm12CXyGHUFnTXYV8I7GRSTZeW9efC3CS9YMLUPUyH70mxD84FpioRice+nH
iZUs1ULPTHzlM6F+Tv1gvU90uANZUL525GEsuVzYVswrWaf23LJ1Ohzs07vvcU3mFTjrNv1Sad2G
pG5f1+nsglO3VBrySld6cjjNPJcMiJO/zLko2dDXoTVxjfBXycjoQbngL6ZVuZW7sfBfCw4+s0MJ
c3iG4bsv+3kZClRa+RsM5a7hYCDbJGh6awSCuBmUT3zTzauDeJLJDxjjz4m/XAJ5Du5yXGiuUyOF
RJ893J3qG7zH2Xr7XbnP92OrtJ4leOabD6d66mICZ4rkUahQ17dD4wRXYjPRkzK2MsgOTgSCLmWi
67Y6nTIBwApoCBBi3pO3EaK9MlXHdwWboecK/ZBw038o7UNSPWA/zgItKLmPCbPmGYgwH7DP9zQd
uGGXuMIGGU4D7I8XZ1da4JNjbqJ1EJfiiDP2PIFRsRD7SMH3UdApeONeHYCTDKLCOCSuV7mttn8t
ToK8U67BrlRb8bNhEwTRJwSuHitQqztodKKkrFH6cDHlCsIP/Vx2bzMQFbOGr4aIHmszfh+IITEZ
HsFGbPE29QQRU5cXbW2dxSAYTda4x5VxI1CWUTmcNdmDhP2Mmzl/dwcFSTXku2phkK9izh20p2q3
Z92KAkRwhHfwYCkkuyQdZnbEy72yq9doUEHglJvEZoJxFTux7nLVeNAOqHRH+kDZ7vw5EF5iJaDn
fROMMO5pDWQBzdFP1c2LHE8Wl05pTQtcZWd6Ed8la1wdEOXaN77kv6K6iih9AjF+rrGes3iFyoHn
lzzjUFlDVjiHhcEirKXeRJcEmIXn3TUnIbD2YBlMDm6yfvSTpLqTRF1I7IXb2c48PVAXOZ5UaOv+
FqIRgSQsguBIWAGVK0iS4JA//G9pGH9iNQGlyKxh14HzsvIVrL6zoYblKcSGRHUNg4uT96d1rZ19
u64KYy5u6VHc69oD8+JMqG4f4XT8GHUXjtRrYaEEwUdYcsyV7R7fU8JqMBnEot9KMvsewXVVhsWS
JB4p32n31mrFXSu9DffuM9HkrWG5gDFjULpRSS/PA4Qbyl41Pse2JqIsNDoEHjZYXPAvtu5wST6j
FTLNr0tVB078J7Q8wuwjV+Ak/nCJPdxbT58kS7YcDBw2eF/uoBM4dP/eYx0yzLyEu9JzdmCH400o
o7Tsnz+FB9l24Kju95JRF+wkqmT3GDeviYZPWkZBNzrsra0x+ATPjlipSi+r5fZNSk7OQEyD0BNE
6xs73gOeCmwD4Qui5MJwUlB/35nM6XqlQEvbMHRpbzENNRSA5qsly6OkqzibAM3ST4jsGz72sYs9
a8xDRmh7oy26N38UpXjmP8E2qxqKDGjqeIosdoj9nF0x9jbuUQxp27Q435pkaW8FblO6HfgBPIhl
b2yuksPrWJK/TaPK/kMUg2KseKpb7NNt9te3lXveTqwyos3RqcAjyhiSnH6/qk9mSOi8jR0DXwmZ
rYZWkF6OpyCsuTJsqh7UD8DCAPK0Wc/vA1BJ8bnbLSZpsdhIvfJKupiG9aZ5zUcSzjyIuCWgkwR2
U7Egg/mv/SX8Qmz18WjjHFsjGeT7IoTMQut0LhjfLHWmPyowFs4EVLt5tHzN4KdCBgiWuPqELpm9
EvXl4o+JdhODc4nCs63ZSJOCRgPkCZQA/mO95dmPXnRIjUaGzEZQlhBtg6aJ2eLsM4dXVGy65V9V
/R0EzZFDzUe6fi3/E4BqyPG6D18jar3/yOsvRcyayMyo++GSFC2DmZg6tMNYcAkWD+dYY0ZdZFhO
58+obJXqiCfAJGuNb71QCb36rpzS2lw96A6CEwxAvmdohC7fTxs3EA7x/lDQbX5Gve2YxLAC0G4k
uv+pQfDAJsRaht7BkC5cYuNt5olK6gp4vEnGPRWM1AYMXoHNPOD0lbCrjC5OnSA8nO0ywXz8ldyw
65wkN7bk4W98cGMZp927QdTpPcyG4Vd8zo4ketYLoSDY6rYi0veGoesB603/zgBdG2Dmv+jLXAJe
7+Ih/Jh0wDGTB2MoJq0OF88pxAYmotXlZc23U5KL5Xs4cJ2qFGTa7AKQ2ZvPqk+xGTyyO0Qt/RHb
i0t5VWYnFDssedDHG3cUiTm3UgDpqz7kP7pMuoa2FsZ/MWz7JDBFxHcO/gmOmHzV9gMjnMfVu2b2
06Gx4xKhLRymHPr5NeFvCzma5ze8/sG50unw6bMxUCx6Hzgd5vPl9x0lVEcJe+qWg2cHFhFtjqT8
bflHXyBS78wVdIkdfB38h/g6yWmC+3jIiwIQnwdlXDeXJ5zhgcyg+SFrFAqzZpVEnNnGg7kH0zfg
KnZOgOLwB6H38xD7jeGchRQ3mNj8BeKM8PTUXP++iB2is6nddCmqp5tLuaA6kWBsL6IHVRcOb5Nc
IneaCjBAIf/RLZR0tAJV+zPe6SLRIOME4QfKTs9d3ybQf4ErvIezGlLa9SQfW8j2TJVcyJcGkbl/
/HjdbqgQ9uZUZapltwZQtDSf6OZPUBj7E7MXqzMVvoa9KZWJk4Sk6qpYdgn8Fr3KA0orgod8YEdQ
E8lmeIKig3ViKOnusxgYIaG+cV/AeM4uohkCUiOFKgFTa1PmPEYrUZfMIk0uHbUU+PypX4abEvvP
z29EVu2TEAW2LHm+2yK68EQ6OqdixIXwXKH5xmRf//Aq1vnuxaHrOvj+Nu+T6crnxuuOOFxQ220K
WQ+KtczvVxFTLg5Jccg1zmDDpOEYf3pwDOaIlULTuDXyMa4PqkndsH3nTCv0lTrT5EgjJVYSYVEi
o20CzYfe4sw6zfFy8g2oUXW5GWaWCnSVXqtXImmQyT/ybdRIxC752tPrqgEIaas4VW6CHKRmlV/1
jSNfEVkkz0rFW59+DAprpwUbnfqwam6xnpts7/NUZhjAfkdzL1MWBAryF/NGeFnMgeaG2Ed6pAZf
J8Jd3rYWhp+FcKdnll8hTDjzeFGOtWAOp8OcL7tMeCB/hs15qaxf38KgWKKfRYLZUgs4er+tw0tE
j0s5dMe5p0yRGahFYNC6Eyk4XEFK7vIk4c8egq92/GCyRfb9vigqeUdD3P1G6v4e2i5FhCAQfQS4
nYF7awRUQn08UuA6gaEtoXJbAMuEwo1CPJbli3Nz2Uonc5GeizU8POHr2Dv2gz3dD9jeeCDKUNRS
Lp/GMFw1BwKVkGWRU+WpiVGMRm2TtIZL0eNaIqA8zitRYOv6Zxp9sbf/i7jKy8kn8SDO6OGbXihH
3zdwnwrAZ1kukbhWl2duRzcqJW0xL1c7k5SLOtDKmTPqducZzw+EILYAzAHoJvQG2wP1dNycM+xA
BOZb7O4SZEWRguHoV5MLL8Bs5iQ4eaIKbFRk5tDZNyF5Al3Gmikn5nZ5ymquF64jT004BfWe541G
EkS+TPAgmR5fia5wGdQcqAuMMJYyotx7zBcO1Z/RsFC7RgXv+DiQwRLUe0V3WZIv5iADuF7o7c06
C5GzuI3OOh1wOa87jOfwSB9jw0kf4KsTX57HH3jKClhmMyUvXs535BUSTa7fS9TgUkKdIotUN0ey
YIUj/yai6fdmWXyw8qiDaF6JO36+OsuTbp2mfQ2g7ODJW/P61BcNgdoVgUul1/MOh9A17uDBvlxF
vDbTJ3FBjwrk9sifjZkDGwNlwPnMnD8nZqim5QL5hlsUQskPm7XfAo1SMDAJp2fpkbyk2QjY55kn
yB6En1oTk7PzlgZ4uoHxkCjXvGwPwuMSOQKGVMhAmzCNT3Er5rmnsKBPitszItZTY1suOmzsHPPm
DPmGH5NtGe/KvN7hJIBmLs6mijgOCHrvrUof/ftd6SkdE0ZcxU/xziqQFGwXazhuJTT8hlEbsHME
2JPMfOCGGccbSFjMzRelWUqx5C29UYD5zQX0omdCz+9UU+JcmM/wdqvwh0NdNGuDtEjxMyHOW7Jk
LabDpzgumOffBup9Yg837Rcz342J842j4mqNThyVXRszY4unOhqCgzrKMbn43thHAXavSHcwkLEp
od1STFR9nj6f/uXWetQ2sAyPmF5YhHtLiVP5gE7+G/EDndUmewWFMy1OZUxD+Z9uoLb4auc9vdLb
MYaU2XU3Slcs7Luj/X55sODceWSWHm1HPrJWI+2yYBqrHsl2cMWGLSS9D3AaN5slAlOeSfnlNYK6
56YRwTzaMQuSJvQTW8HfjZOFt/fuIA4OjEASHEcO/Cpxo4f66OZR9uHZrhAg9PhK4EVhSMJnC25C
2U1rcptdVqaBDHNZ8kryV8uXAyb9n0aCwCI2qfVPsi8Iennrxw3JzANBq8NFNPuKA0lG4XqAwajP
En/Au/qjOdbz73X7soYVTkiH2ir/L6Tk+qIAt/GGJvfvEQTO+coG1N/657JZRk2SPlBW4xTmUSGx
07YU/UDauk97IAqJc5gfnfuU1oWZZiSxicxcgywhWhmw+yptfJzU2yfCEIoN0xWhS8DGy5ZG2mCp
dv9nxeTvWZLTcqrPHzy1Jfcn/2Z8/X2Las5RntTFPq3ZemV7GGn3S4OheDNSizrydPWAYIAessVW
CYwYY9BQY0wRcaQrCnqx328wva6esofZfVTVxpdCsg+2vqW72HcIOFglfmbfh9TKJOF6PDG6eVw5
Bc6tEOhAoT+uq+IVTgOVuhdxMd70QbZ4s5L+Nv3YX4AQAYhSzc3J2K/yMMiHiZrKtMK1rlvNoEcS
jrpT0dpRokWHu14c+lPXMMwSQ4TJnnP4PilKbcCpessphYN1bek8kGPbLggYN6i+KXRPsO+8F1Bh
BHNSYUzhzkFQOnQs8nQcKbtXqTdm33YG9naoswD5q+ydHwtkzHtMlD9rvEUUkwaW97AFOAK9gDBO
JRo7AhQYrWCSnbbPkHPWy1QGi9BHwqbRm87wjNAIrHSUXJ8kgrfYIHdSfsnxy+0bS8ZnBZfcFztb
AmmT9nVj4p7y6rehsDfHI8sqMV+XnH2FdPw3oxvDq6tTcwgtscAtptCsZ4STrfN07n5a41haSuLl
obWNP6ei/BxSs+KBHFkQX8VVTtDLuC8dNBGbFPq2wgtGvFP/G79ieS8oVyEIS2LmqTYYendgqjHr
0cBT6mR7yVw/6vTMPzBIr0Y0qnBY23qvM5RH18cT63nAs6Yz/WrQfvZooVpWVrjllNrjC3oC54tP
hlYtGz/HVjIGrldnMEDNM4dBovpexNnmIVrgtbOFjA+KLsIM/thGvWNHpZN+z+kteZCG9vgi6OPR
g8xUlvu3clQZ3MUb8JonOM9VkGo9XdC9RhPj7MMfRqVERBpSASWja/yLqhoZxWTrs+1m+Ngn0EIb
7O6enuzzhvmAzmsOG9mIDr4ib+zTrmi2a+ry2Q/GKZ6ZJbruPcQxxOCiGTXvOYrl5Zr7lU91mcUs
f8bwL2nhEHRSWmwTU3iDE9QQtRQTb381Kq4N7M779aRUQ6E/FZ1TMjj4FSn1/T5GE+HVH4Tb+pCG
UTHW5aAN7nCe5TtKUoTrGCmdQmQeCh00iET2lxCXIaEIiM344vSMTYBueUO0KP7aBa2j0xLco4Pm
sB4gguGAjepuUCG/R0dpW6JxiOrEBRkCdTlDS4ORa/pwnAuGlDUDs8LfDLlrSpr8bfwo4eWzGdFK
9VWOHg9obWkKpM1vwZoVezYeMgthTyfyYADA7QZiZa3y9fHe1fIMexpsXAUsAUc+Z4oRcj2T+edi
3DGEMpw9Bq/4oEXyW3p5T5wvwsTsv/tlCJFtpyQJQgZfLSjK6AXlazNkY2raRAxvOSpHLNBir7ny
6TLB02y2S+1UKWx0ouwyBZuTWSyT6OGHWKnsFaEAadbhy2ZO8R5cn1SylufB1n+vBCv5UaJ16IPc
rl2afbTqMeica3ByFkEjzvkzJ6e4UDQ1BJr7R5aRV2F/Ng0JwJlmuACGPBVHzliT7DHRZ0M1UGsQ
ypl6UqiDKpP1GTYXTevfcuvuZIYLh8Cbgv4ibwHKsy+Hma8b3cGhzU5dpRp9nn1d61Nbk8yHBkrN
VgsklL7etwJ9MSfVFQaJNbCXj00Fo8AVYc8V4OBgMcFOMPm8f3gvOuPN+oiVbBW1U/HQgbcOwICQ
CvNu+T8wezbv6JnJNoyUtlksNQpfDlGilwWP0+Lu3RkAWDQUohtb7SWh1u3b2DWLbGsl+a6PTI5k
mAnPxFht1ZEGdga/Ec1MWZJ3UyrQy909Fuz6sXjoHwJFS9OwkSVQniP5ebIOVB0NXaLJn7cBNF45
Osrn+bzMj6nnhloL+Ix9oUIsiQS126FRmgE0YiNT3gjEl+vQM3JHnesjccu40P+Gh5VUTijUdl6S
y1RzNLFLUiPn6Zuc11vEQ+wXstgyQPLQyUXqlIVaAdCtmwDzBQnILocViSozyOmCoST06QtgXu03
axaw61ywrdEJDnZgJhDiuC+K3Q2oCXK8Ihr0PCeGX/Zy0LdhMZwyDoGcDN+yOOJmudV4Ylc1M2nr
si3ZSxs33XfNqbbjHpnPfUe6QU1Ait1QXtmcKZBB7X1rkVtttnDUQvHz+iOFykLxLOUHN3+8pSI9
mvaVgvXlcxjzORx6zlLMBK8B+0CzELUl4w41jWJomCUIfug/IvWN22AbU13iOeAhXYeTnob4Cbkw
SsDFsuAL0vMgD66YkpTzIYdAAwbhicDYdl18hc+dpQe/h4ZEgZyW12omfTMIrA+WwL+NzpC3Ii3z
yebEkZvU/PLoE4BqO0JT+tssEZhXAtKMhCTThy54gQzI7NKhmxkXoarS3Wt8PgN3Si5qRI1GjTbr
A/ZMc1fpxdJ7NWQ3ZXbv6Wv3irAVWoFXR3CXG7/qLlFjrv/xLt9jopVkhDbocJaXUe+0qO+AfVz5
vC2lTB55PJ2f7/iCLX9ASDr6OA3AwnlHJiDcrRQugC2i7YFTg9wbnXSR7BnqZbqTYkh7Femf4Jxw
4Uk8FfY+m8l30pGFV7axM6aIaYyfsoXYrCi2vfcbvagCcoTxygWM9cmNM5F0Y3Son7kDTmC7vMDn
RPitaaACSoiTXw5h1gI4fapwoOehb1q9LsPtTGkTN5eA7KXZbyqXhuLKuylqxJBqFTq8G9/8asXs
H+ZfUqA55Stc3gtsLooAGPSGeteBEx1iiZQYk23adzjL2gipqnmyA4IA9xWSWnMIqCL4XQZVZMQE
9fd9a4ot56vEt7hVkwdeCThCL1UCcCUrPuWA3YavLDGuDcnagRZW0mUXda01HE0LhEk8fE78NAGS
z7YerIMmOsK8VOTlZxVDH3FIX6bwNUBp4lOYVNIyfdCBGz/EmUgM/gJ/Tzf+Mjfy+iD5LlvFaggC
I2fmnVDiPsOQ96HWizZCQpoO42EFwE845eZrsOAkP3fIR4jqhfKycdTu+u7bEZW/6l0YsXE4oW0z
4myVqr1KbZ9gdlt0B1iwIfNhXKETw+b5t8/VYO81sxT7QzAN/s1v85n6OTtwtFi8rqlt9xqkcvzx
2GnPyvwroWyJwmOYVJPfnJFGC1koLH9hu3Jga9/mVKbnR9GNuyOqTd9Wj5WVDeUW/aqAqhsTYpVb
jx9D4EAemWKWrKS1xDStX8e4hecHFcZc2GTSrAka+wXXkXkuR0omEHCcdPDdnz5H5+8/jRnvb7B/
vcw1tvBMFUDjmkZ7WUZsYqikIVSKOaK5CT9J7U17wSgKxzQYcUsjL2LWyp+DEaPLF+mDzs1KcYlh
ws3yKLj8BAfYX4g2g05a2jDiPvtWEOisT04cdjWyNIcWBZXDIUiqKGkglHBeFhnjamQyQ4JYUoEI
y7AwX2VNjwbBS59/LNru9201Xio9fevVdLHZ7xLkv57MN8exEeolvDi+vvrdOcvHdrPqOFitbZdU
cXth4up56rpcbm1lJy03kuTBAaGAJ8l/Jde4ynP3EHMCdj/r0roIBefD2UWN8311e/IPEVe0db+Y
1Xa6qZJAO8xcLVmOvNArPzH9azsDAiXbFxb98XXFTdNPUOb1KclFnBj1InoaCqpwYIPSmTh0TuxM
eCfwvDYQc4nQEqugU4HsLq9aVYNU7wpq/Wsj8WMY7JjJ2LcV6mJT98K7TErriThdPb70mBBVmOHC
5V+PPIZFM9pRcX4j4furGbTa5yBGDfqooXQXAuFNdMFgVv3j4O894Z5/Gp4DpNRpEpk2RJQqvfAu
vcMqlx4sopqFb2LlVL9OQrm97knOeCBgUrmC8zJ8ZiJSh0h2Zhjfw287G6G4bL6JKx84mp+5pmSA
31qRKwg7hQWF5RF9bjqZWQgan3Nwvd+KnS892Gb/76IAKkUJWwJTKsZrYGnpYb5AXpp9nun0ggiO
QTZtZmuoDSrRONPauBIlbo66fjJdJ8N3gvdl1LLhvkuvrdVcz5UKjCgkZvqq7qgIp1AoNeQpqOh1
Zk3Qmidtrzp/EcGnkJ5Yankc9v/AORSWWwVYYEffqSQ/tRGuFyunK6eZa707cbLpdHOauPQH52dG
52epN/npwYGQYj5uZC7fTbeCHpH8CKXDIJiR4Hr0c8lo2J+q6Ckn6YHYdSo2xEDV0/gftLwirJX7
EKz5/Fyub2QqhdbWfAaHZcETu6tIrag71PSlCiEOQlklD9Shd3C0Pz1YaPv//XU6cA5ponx9frDC
WxtXDzw4kb4Wj87GWXdsbZJwf9gRYIotE097qaayU1VPXFUKzH5eGrxQQEcE0QSQ27Ff/KOGmDFO
883pbbfQdE9SiOo1r9tlsoRbGjfegEF4x+egY76DZwbgvniJqy6rvgm0EsA9YWpfCv/6JaPJw+fL
VUdKFmVZfc3EASP7aLfxtAFBtm23GOTaT+W5tMhUzIRC5KfJJSTosDYWAgI/V67z259ZVBixlEBY
iwg8vu8ral8+VdYWUYzB2qbFO9NwYQQ4vYV10ZVx73+myGq0sqf48trKHE9AHAxzyqAZNC6I3MpV
ZGd5WBsvo5vlIkFYn+TZmCAkCD51AJJj5K/pXtK4UURVAfKEBy/Z4YSCo4cqy9/ZrOCmYWXMvhlK
4HmzYyvSp3fr1UT5KqsqY2e4LMZgpK63I03HSh8n0aveJ9OZSHSa1w7H4nmiRmdTZotDhjBp7fi4
R6QwaYwXwYIqQrseH5z2v0U44DZJ9eKa3xAbV2M4M9q5laNLwvbry5gGgC1eXtPlvP0fj/xKjuZu
QVGmJl0qXOhWLihxwx73Gh65EFSGzLZ6UaRt618rHA50xzc2CbhvFVGZrEAh9WMrqYCtJNgIiFdf
ZmtX5Ey5qS1m3ck9kalH3UCifNek4xxK2EUc5KVGtGkOBz4lu3c4C767teCDsE/4WDcMlOTY4KJn
/HJ5Mejf8fKRbPh3JVVwpbVA9IW9BEijOjeMYLbIPPzhsWgRYKO7jHfEX8aaIIXLz6AvXzmINYVM
wRfjHs5CLDnuhi5MO1/VKA3yDZ4P0bLXv2jGfvGf9nnzCGBmv0UKlpCcSjjYBY9jnSawNVMHKS8r
STg9zJFpEuC/kyK2TeqjsMA0atNhb2yWKgThbOazPI+2c39fQUa8Lj9m/Vbn03ofkjO0FJfvpF8c
DkHstW15NZPTnBDgJiwiXjHlFxPFsftGnpvsWb4GW+sAWvlPXLiLt4Ofrvc3mzCyLFj75JTadi4s
94n6zSdmF6K1IyU5/kFiHgDtG22u6AmDJYoM7UG8XU8y29ZHqQqUJC8XBqmBbg+ybz8nmkA34cK/
xCCmmz44S0WWV0y3EcPyYm+aS7qe3fwn0Ce4zcIbmOUPSUnYaOMKKb2F5vjzl29WczPUgnn7ImIS
hb5U0tv8RLJocAMzn0Zgzz7AzQZ48vfqnBgL0f4x5tUmQgj0hIIUxZEuTVbig44RRJJUGQ+IO39t
weUUvxO7XrPB6FLBbtBIj/XgwmfzbHkKgjg7RZMy8ZTCtPC11aWU67tYI+YaUf4fIaUHERGGJ5jh
1sAxP9VkntEzHzq+QSHWx69y1Z9IoanhHCiq8BFkgMn5LGOXTFxiA/urQ2hfPdWk/ICUEmKqixKb
6Y8McJHhGeKZLW4s7pQB8j54p3OBBldWh/ywoTliwMYQ+UDxWfbQN+WK5GWsmoEsxXPAniZiDZjl
HMUloBmD6um1F4T+xFWDCE+XF9pIwL9jZdgo0VSONh81hI7fav0bPrNqgyIjg8HYqlXvHTgxSCB4
HHjWvHqQ1GP8hz+ZvNP4qnVLhLhLtxOdcFytEFBZ7sRdmNCVPbFzqyOY1HlPfEGKbpnqsQ523Wjx
LdG3g0LPbqY2TOkNIlWlGilsnLGBhwQB/rRNyDomdU4/b15nO0TrHIpUGrDlkSD+X5K7rH0hYkfV
ht8xCw6iXSvnGpF3ln3cvX9/1CmeG8d6Y/E6Zh1BGqrJMrBC5BxoqETXYqDmMd+916ON0q6q1E5F
qXR8UiwpsiyzNNzIoEyjnwfStb1sZrwN8kZd48fpcVFf9p+EvNLBaTCJn0bzZGEc9xfsIGUVqe0o
t1cdYUp8Jffe7p4jOmmuE2yozsshLyyPn3meN/fQM62Ewnr/qMI1mYRkq9sMSJfwtS0CHyDnUdKI
m+DSssA7pKEEXPNf4Lkb5gwenZcDtx8Ot4mUxlCPkW8ra03GBcNnQK/94s5EdAxSxbtKDLCrvWfk
qPZMvdMPFQ05lAQGJm4QVNWmEEfJX+ovILEOdVWg2enU87+WrgWDYlMUvMBXbPgiJfN0ncsjJ7Ss
kaN+32t+2LxP1klXjYrwCC1LwT0K5JDymv7ERq/00cE88H2LSPnbZqLoA7OGRP8Nm0Vwx63Mcliy
ealDshR9q9JtSlXnbV83wDKGDZPx8A3N+KiGtWq60OnycoFnZzgGZfsxlTddva3i9+zyb3ch9ITM
kYk60z+g3UGfjJMZySlwbMAdV72VODOfcXXeOtOYuxWUjhDCD4r96DPahX96c6CNMJJh3Tgv7d1L
QFaxPD+drmG1NLPxIhDoH1ldhF3krC/oiMtLGVzchTo/ZMj3rVOZhJIEcobJpBJbdxqYbKNUbCmM
Z0KhK40niP4q/dgDkGI3k8DBigytbgV4HVYrBurGpaVKVEftqpk3U6NNjdBtdpsw93AZklt9lUkI
ti6+bIXyUvD+j+yd+Ox15hxT1FiNczJHDEXD5qCuVYUODkl0IWOZWYjA4v0tdLeTWPV8cAB6qaZ3
tUoL1QEUSW/5dTzr1EatVd3GtIgbQDsoYgTqdn/AS4Lnln0vPaYhta9RGk4fXrWwNLyN47QZfyWc
X1emfnp2ht/SuycGm4igUBIiu7j69ZMhiRoa75gaE/nUBeZu9mbE8KgsVVSThP8qzenk73rY2auG
IG62Wqa/Pd8MDP42zFLqT7deDnwmQUVkVYT2fCXhqcpZExZuyulFSUqZ6UpILwou6ZuRSZEX4tCJ
gLKv4yA/DbTz6kfthCcofcrtKGMmB+GIqBXSe0WJ7lrQrAWlQpzz0Yhn6jzWCpdZIEAOdLxYNZkp
/wyA1XfsQDozeXPazNMWbtPlF/qJvZIklB2gKAAjXlcef/ph/V9aUb9j9dDI33G2Q6+mMRn6mjXw
UvFn4Qu1kFr6Um9jWrr6RnlKWn2PpRXiSZt/E0pCcmN9HmYM2CfVjwi4GhvSh/ImSUfZEeMo6TmL
9pfEu3zcfPfgiY5ioeEcuUAq4IggApW7TmVdsEqCD4RIREVJLaJXXiHsdICMXTg+JxaaphrPl8l9
6mM0mz6i++NMb1qN2F2/+VmBMCClQcdppDAE3Uq3GbIASfXM7U0w0v5aFkYjrJeVs/oGRv+k1c+X
bMTId8cTx2QcsOBAlvq+6PgmOIRnLpv6d7X0Z6JY/Yhm5JXEE/HdZ6xWRzz7KU8jxKIh6gNkQso3
9487WLwp+zHvmo8bsZuIbqvAPvRGHIxBFkgzg+Gk57VrRvdfnpxvAEk16duf112EjohUuUrJtLJc
Jm7TSNlKsdNM8kLttGXat7V2Ca+D16ftfm5caXBUyaZ3lloqy+JmTHUiLbfiQloRTIcoiN1tg798
fE7aprY9j6IOKLb2kE1RsGohPe9Yf7nDjjwjiAZGkZjSX2KGKSyT6XSVS/88G1pYqeNeb8Atiz1w
RCoYTT7gItcF6XgLc11nZ4LTqfa7OOfkCjmf2O4s/2OYqSdXntVM1ZT+udHlDsy63/WkVKSxw8e2
6s0ESoegMq+yDppjs+F+OjkvFxPfZO6wjTzj0nC6iFphG08xiGimfCget+xBSiFZq1LB7mVtyd1x
GPGGCo1x/9GB9l9QNyLdDkWg5abhgk5IMLVW3vC5ZscNTe8SveHFwS3IunBwEJG94a0fzIP+cCfp
R4ajgq54+DQBZeRmPXbxh79kDNcwXkHssyF3nyu6v2cCMeCFFJob4WBEWyyAom2aD1PX6D107Nmh
Bxkq3chYPgURWfVoVpJi8i/vB5yiwraZq81Vs3qgFy4abEmMWs305BM96cKnPq3WKLlZJME2NhRO
c6vkzs3xxSnMfjuRz+LNydCfgfvgMdMomEJsfnBqJVcNNHVxr1fwsk5oH9KJf4/aOOGkzqEFkW6D
h9vwGWbDwJW7rZBzb5LRrPwEBWp6YgRwLAPF8vbojpPLEoEXhcx5aW6LcCZNEgKC3F5lOjlgniaB
q6xJ2ixYDheBB9MaWWE3YIOcQMJL4I1potZCRPJXsrg+Y2dlE5IugIQDTBV6xK3XMflrQbUn6EkB
Fqq9JABj0qSv+xqdXx4cwZe45my+fO8r480B3T5sVycGve+whQ+JS19xMkACKQGdgNAYzEH5qc1M
pAu1tJ9PU+/0yFE/yw++4duzxhP+U1RJ+Pu9vin+C21UWQ4QHsuin5DctfYBkql3EJz6SP24dOJ7
pg3p6C2eF/+/pIHzw2h0FKtoSReCCrrsMfHp0SRPxpm2gxDglsJQs+zoamGdgxF3/M+rbcpOFeUu
6wUonnMdTyA7nfgIie5EQyO2AZXeUR0DuDILhj/XByaQbECZ02ZdimugEGA+WN8454F32BBr6Gtj
S5q9vqvkSk4EmH69fm4btCLq3bJaF4+JSbrmuKUWspkoz++OZE2n7En72P5Wv+y8GE73oJy32KLf
o1ov9ImI05xz+q56z6gbaDuUhzz5zsJFgGe03XbD6LV5+rI7M3/LyLMdIZiLmL8pIFhGCXM6OjCQ
/txc25kKUzMJnq2/gqYh4EZg3sG2dtSWF79g/62AadCqo26M3+h2B9xSncZ4lCP5ZZ1fIsfuYBfM
HRIvTdhToYETDP08ra23bu06na+dWeqgYeuLIo6ZVOhUdi9WFjCVgZuMnj3Nangqzjxruxkx0zu4
6Elp/IK9We8HkGt84MKrpTQBoPCOqlWnr/2xLF6/DFzfEV3N4ULsWwwEuUoadErvrY22O5KO9D+8
3mSmedbZtOQLmxPEaPiypozRST3viX8/Bl/e50aMXbT7aKt7ozSN95UO/y1IGFIBsWAIHqi28BuC
vYSxENjK58S62mD00ryOyDt1BVmGnTZQ0w70SqVnM8Py4YDp0cWeBDn9tyJKSH/gnxDJg43E1Ivg
ScV3/zWOXLf+82+wKKvteR4Wr5Jrf7x0+kNXaIkuuS9a9QVdrpqon2DmpgJlVTMltiQNZET1ZrwT
vaM1zVOtV98arDLffYnHpBvtWPu6lyoQUonA5hIVsri1/yO1v1w78swKUM+GmW6DEhGU2N3LTOiW
U2/rrtZLjC5GaeCfZYd4qwABijHkTgxuMwRHV2JgSbODEHlpSg2jZ6PrmBNLzvdtj8vrfkECuJ9E
k9M7GLbyBBpYRfO+qH/qO2jjv8/WDj64hHSc0DNrTN8q+HexaGgMjSAKqEYfy0hsFfSUukgZVkWR
EGk8HqZpPlTr3NHYBO+QvLlfKQgPspRl6LepuNZ8a7E8bNxi21dCghPpFZVxrIw7ryzb7fT9G1Y1
ielbpI8WSmlDBeiDBhT4HGeZMCB7IIFnX9HySqXLIv/EGrGNBGvxL8938BdcCP5/1GNBu5pm90XS
TCCnn/uj95Y4avVMe/+OvLJcZpQ/f1ufN6Eh1vAQdp63BQeOvToMrZ2JCr9nCLOW1DJ+hOXTI2qD
Jg9MVyL/Fzygnc2uXG6lGAxssunhninjrLE/cPy/3P3hXH44vuVUKB+OMvCEXNQ/ZJTMZ9WArcvL
73KodackM1RKS8Jo5Yn9EyNR+oimPCt14e9bpsatXglbUU8jzkF4C8/tIDuDlrJ52N4jzi3Utd4T
W71yagINVDJ8Xf6QEOXlHjiUj2Jo3XwrCbOMtk5MhhVuUepuq1v+wWUJrDgl0G+bE23R0c27Eixw
Zzy6WXvIjpkQJQS57zXvUdRc5WQnTALrMmS6qOoT8isPboHLVbfXfztWSYlzy+nEVa/sFC0Ze/v1
RbEF0Tn1tYtbE+wT1lP7xdZTHXwIuzEuKoFq1ACKXCjnH9vE6wD0FIpT1IP+qlmSIHIKknrONn4a
+gaJyv56Vh9Uexu8mcUcaOcHvntXF6P+ZTqKgreBjfwTb0qeaaGunnbCI99Wwav+e4ldEZKnkohA
kFpbxh/qMXEf5TwDQ5i4+pvbRUERpcGny4ns12zRu2xcE5KxtV+d6IaviZoqacObo4Tw0UMALLOW
DRSbl+i9/hqtap/nN/wz2u1NMgUcICWw520ZjMOVbSMKzKuq+/snxVVV4yhRZoSwlJX+b4UeQL9E
Pl73+RecKxhVP+v/rj/JviYA0oofhIDdEvaVvs4lqruVutNcpek5TjQyGYlt6gZXuFFgcZGX2ysG
rD/6sUd6g7pzviIKq+MeKgQYLNI7Lc2TZu2txOh1Z1sT7Ga25v07YCVwzpkVMlFrToTiayo6L7K5
R9xyBevONdjusG330KbgKkfQ/8fQbsqqZGY9BjDg+eN5bONdIi8augeFXzKzgMO31ilGQH2pPyOV
q87lNRed+0B5onPCAyNFdtq+aqTyYXQRDPzgiDx58FMRr2wVWmtdKyJA72iucmaVnSjTF8dZh0a1
z5EY/zeBsu4ceS1a3wSenwxFhcrwI6XYKCRpZztq81RdklYpmY19PrVYWemh2vuE4ZC+pAE/Msng
I4r0xHYJ/7UHUXLRAsYP/+rHtIeNFIo1gQHOkYHlcIeJn4C5xQh6DDACpwNjB/9vMkqzpgPEImQR
DSOMWNSWtbcgygp+lsKaKmdq/83vIAnN9KYfbuWPYvpTNMv96j5hMRS3300HYpjXEzgEjNpZfEXH
qYleXDE9j3LcdWTTVscjz1s7CJb7C2tNMY7iWFY4Iyes5IS/2HkLr/kGk4Ae0poUnQegpVtFvICO
Gb5ID16Pv07Wg5yNEKu/9XnkMkWvTHtM1SPeRSADizqgqVKuukcgZ+o9GuIdtr36zPHHzWCkgg9K
lJG/++2icOESMeSRPGpDm9zgsTsxYS1PKGFC/DXhVpzpZPBVhKvOlbzab6FWOfawdovXGhgx1qcY
i9DvKovdI5CWC4eWc73oqCyWYfyKQTQyhNKbAQgLczvAEXRt3hQU6s3hVB7gJ3+Xp8lLFxBtbQuK
ePadehg2Mrgdqz84mZcVEizAwc/UGpV8ZWuakRd+nJJDdXZjCMmq66suR5xBmh5G7wbeoHkkD1yx
oSj9slBf8RTVVfbPbnFucEjJMfWLJ3LVdMZc+1z8LdM2mJmy6Qk1i5Gm1K7CVCyRPzRLzdrRLNPF
ISH0iDGMmZfFdNmnHvNSUlDeeGD2ABvcbfJmHq/v5+x+l+1+/O4iEzFJ/hmFWH7b8QBxBPYZkvOb
RNzjsidZHRxUqnvJer9zr+bxWmAXg+Acd/nERbE9Rp3N0CXHnSM+f/Ks5l3qlyMLKis4r7YS80e6
fhYuOFh0DeH5DLutkMdCQF4zwQPV8i6Mrn3K7/1+dlaqgQSzRT0kR6bUpZoIHNBOOAqi61NXjZpo
I2iw4uCiknGKv5L+gk70PbN3vQePkBavBfoKnJNH3DzGTZ+3BqLs340GG9moLQ3LQHt1VCpXmB5j
MwedMg6/XOtQnc10LSlsFlq5pWSDa1ypndYFrx7lVEbR438YryrnnNq4wQSQPCEq9FglFJJsjkLy
pbRlLRPDQwJgGkf95Dsdlv9NlN50uGt3/PL+7JVwlU265/SMucXkXRg/MrRSDc+HvH8gvETbSTMz
LwicYc2+sm4BHwRKmqnviJeYsObG5Qopg/4D0sumprrItUpT+02h8TaMxHU4ALUTivPtFvx2BR+6
YOqB3Z+NBggo2Wfb8WiNjnZKBEOfYldUs+wO28amHu7BDrn3g7rHs6hSfrTWojglieYjspqJke3A
6wvbirJyvnVaIkf3f+UOuQR4x7JGC/4chX77FINO9DIEJjjTK/9ngZ/OP93t4PX7XxSvzxHY3aoC
i8PrlJc6Wf/6j2yYW74mZGMuCrGB7uLSwYkhhNObU50LCUiIPAJhrCWMKgcNrcky179xWsLOLRcz
5Bs9WPLhbjQtgmlp1BPbJaKz+QRpz+Clt+SSz3FO15lOZpWCz9OzNys8GR+3NvyEclPHQbezJwx7
xe8b1xMYUrxOl5cKFF8KaJNfWj80md67CPd+jwNRu4MScw88PBmCOskTgsmj59tHiyIncC45J+fZ
UI92ACbdHz+YGqaG/gtG3srmFQkyRiT06h9djXqlAJidKSeaaVYWvL0qK9SN0YeP90ngPD+jzibG
KhppcVv0cpWGHVCLp2WzwWeWWx2jJK0DFWjxoCto9i7j6v1ehERaPshxC5B9h2zJMVv26IxMJ2DD
p3Q1XOMqdm241E9MUAkpaEy22cL17MjngFsxw6f1mKX99YL+JkNX1IHD/S9oedwBsvn7J4qPS/M3
DbG6+p1ZxRJVgTwcPyIwl4qp6b1Jwta9Q9mT1YCLBUO5WLzwNtH9acNeMuqCp+AjYIlnIF8VXut/
quDTZZdkZn/jb5pfhPThWeHd53ZWG+pXSdLT18Jsk+bl7kO3cckGc8ROQXBAWOpsl7dtIfrRbCI4
ORZNqtDCBerC7q7Evu82sMUfcHky+SkD2ULRJN/c9mRcGH7fO0V2xftGlGfaWNubygcY5i3e6s3a
M0L+Gh4OxL7r0GDh/UJpTm3+VwPQMOfGuuta5M7TgkCTIvsJnqqVYqnyjk/LI2UV2XuTZdjBK1BL
Ttw/RRBpUiKEkwGPgkgBV2hXx9NnlnDrya9mG/JO0R9KJyGnHrw4bAl5koMpOrGw952pS7+98GnM
UL1CMwpJ67cFKHYlngJr72tDhHW1/Odwj1kG9Z2Rn/fITRVbxoMo9aaB7eSD/jdHRfh+g3L6dKkW
0wwBapJZ7Ex3bb0CSC49dTu/Pky7Ua+SjnOIbwWskbdyUm3K/e0cIJKzz5JDNoDGDxzahmaNp+SA
YF1v/bglXtP6AFSLQloXfu4DrgTm3SfkVZpJ6bl5vyuDn4V8ZHtZkq2YZvIxZLtHxRZaSPNfG0c6
iHRLmOgM43OtRXtlPLh4KXZJ1a/B9nsFcaldVxKk8exTj+mgPiQLbeXV806bNW70MavBcOZQ97+H
nSmlLWF3bhL5C/Z7Wx6O/GxPuiMxezEjl1vvlhfCQOoOu20dwUKIU50NIOJvE27BLAczWsA6rCCj
SxICd4a9xHhGoDkt/9A90Z3T+leK3INU/5K1RLjD9NuUkLOFZHF5oo5ycanLCNZ7zodpMr7IXUOU
gtl0qMdh/Nli/GC3bMgEGVF9QJFG0BjilWLPgEJh5v4zj/IPx5HMIitdl1vaGRxw+PyfoJ1HJMrz
KoWeprrlZt2/D80Fv2Nm38JC/VwNR/soYu1uiogDoQOThzOw6+HyfpUKyniI9afrhAfjl4SafvkP
9fy+/NN7zf7JuYQLRhTH9bianRbBsuGJa2C1WKFvuVGqy4XtM4mVGDcsgubjRk+9YvRcoW32UiKX
U7G4urnya4w26VVUFStK5Az7Z6V81qzTmOuVE+LCIYQuq80j
`protect end_protected
