��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����N~@#�k�0!����+��=L���0�ԴZ�2�Mc���ZO�����=�����վ�	"cqw��a��TS[��{=:�����K��-�մ�(��k��N�-� 偙O��QZ��~rL'�x[�i,mׇp���O�I43��4d�,�H�����SN��d���3���r��m���̨T�I;uj2Y� Er�*p�Q$Gm���p�V�`�2^���,hz�<p��l�Bxt�5��s��\yq���#�@W���f:m��T�	,*�񞭋����_��㧋l�	�\�:��uGd��PǷ��N�I��_����Tuv� ���us�(H�~�{2H�:Zor�Q	#%�3ˠ!��iS��95�,?�.���/�F�i{#���Tp5����Ҥ0{%���2vpn���X�����@l����3dc�ק�3	�Ed&3�ZN O���z��s�yxӡt��v*}ԫy nj#��lc��m戭k[��5)�A#�����8�!�]�Z�s�M���t��w�!��'ÒE�rv��Ϝ�c@<U��\tq+��&|�&X1)C�����r�A~��B�&�����s�:n{p��͠R�X⺂L^��R����c���f��J^?��ܣR�O 1�rV���:��T�4���AD����˩�F�w��)Dm�O�b,�a���1$��c��7t[i2>�ޔ0,S���󧇳Ϟ�ᒨ�-��}�!6��Jyv�醊�^_�(�H�(y^����o#����X��3-�k\8�M�T�"`R�DF6ȕ� �,5�;Ҭ C�k���1\������k�t־9�}���� ���QHF��"��t�9 ?��{E_�7��!����]k�j*�Q��~�=�0z����o<���_TC?�];iW��M������O���R�$�lIlqֿT����N�B���ڊΑ��R���s5��yEK@aTaz�]���@���I(��udz�Ȩ�k4�kW��Z�����ؼ����cҖ+��l+4_�*:^*��-�����IHXR(	�҄��e�X��܄2?iUrcᓨ���ً*f���h2\ܲߔ܂��2����&n���H`a����pp��z��5Q�`�sXn���M��l���B|������B����"� ����3¥ ��g����?Z��o�w�ȼ�ZV�%�������v4�-�0�t��}���`��wXXv߾>��%�6�N��_����d�&w��)�+�ښ�]÷V�䵙d"�0�CB!�E���l�Fr�gSaw>�qE��}wJX�򑎣����}BM`\qU���'=�ww�@��],�iYd�-m�M�X7t��M��o��|��֠o������UX��ި�5u��Uŧ����i8M�UŀV����cd��pW�8d6�S/���
��&<�Ջm�O(�t�C���!��q�J^�n�:��*_��Df/�\b�gs�6�ޏ̩m�w
�3�|���q�LyL) f�`�#Q�Z��M���>R�Q���6�V,��Opل-')��I��XհK�h��Pe��r�XO�P����^`��l{B Ώ�@�+���7X��<ue� zMs���Ԍ~��#�<�C��4�"� ����:ш���W��eLV\?����p3�G�:��h5,��*<�	�~3�0�x���ę�������	k�vOZ���={%ʝT���0b���^��"��C$/�Mhz��j-�E0�~�|4�u�]V���;sg�̱�"���pIelA-6�nd�/iHbB}X�h�$oq�7d��gV?�W��*_K��Lh7�-Ë�zi�M��?�B���_��^D�T���E����.+�г�8]��y�J�͞,
�74L�'���M]�B�%�G�������u�wP*����@�w�9���7]�LH�c@x�|m�p��9��}��"�1���=��AT��	2�_a{�Fvޡ���K�)<���& �G���R@�hk��]�VjF�����h��(�Q�YL�G�L@0�g��o�Ļտ'9��oeI�)b�����}�}���·�:�g��c�b�B*�E���L����sS�Ӧd䜔���y�?�#*v����|-H�*B�^^84��0�H1���g�WƱSap����r��Tc!o��(C�<�"��B�Qg�N�F�3���G��%�)sc#�x�B@��2ن���8K/�!�?Z�G�-�5��p��=���9�IK�nEk�����830�wм{m�_��ے��g�V#�f$Ȳ�L�N��t{��9�����c�����=>>��/�kyZ�&v,hfc,���6����5s>xR�|WF�)�9~�
�f�ͺuaZ Uj��1>C��C�I0��1A�j���A���pW��Дjϐ���gҗ�ڐ�n�Ti�	����+���n��S1;&=�����Ұ�Z������me6�`� @p��pA�,nz�y	Lޡ��*�b�Gh��а6�-���I76W��?OA��i�v��H�I�>M���Bz}�p�D)�ֽ�SԲ���W�>�HkՉ��8fN��ү"���D��#'u?�n<��}V�c��<�ʱ�kķ,#j]I�@|af@	Sp_����o/I����$�25��:�\��N5�+�DѕK�}ː�{t�j. r��@e���6B��·�dv�)�E��S��y�dΤ�H���a�b�Q�,���i���[��A��D�Bpd��k]�J*�����!ON��'���R��02;k�uR������x�Y!5��[?�I����'��~��ń�S�p�ֵ\��<��p�L������9�-�
��U��EEA(��cAT ��e�\ ��lHm�S�j��{����C]��GدO�W��������kIg�w&avA0���f��4 ����DT�`�[^�B�U `c}%����4s��6�uv%*u�g��-�(��Ĩ0�.kd�К�PM��N��Z�9��.9p���>��$t�x�@�Z{�
�d�(3}�)��#Z�n�
��E�V_�7��pY�@�ju�KK�ϵ	���3PF�C��q/�&'��HA�|n3����qsjA~kL�j�5i�p�T�_�R���j�W�f��,�.�����.���&3y�=5:��cY��;z�"ɦ��d�j��_k���Z�y�tfY�G���nl4p�N�k�j$' 	F�M-6���=à!b,���:N+�XS�ZTO/���i�͙�Sh8�?�f��m�d�V��������G+	�&J�@>t7���+ M_F7?���t�\u�F�P$n��y+)�{:e���q��XX��I��N���O12LH��� �+����#$�^j{�aTQ6�����WU��I��_Q&�����䵄��������x��}�ۙ��j�i�H��nd���t;�우��mvBoY���⋓�F�噯�+����w�(���#-����g����B����������'���vr ?�hf��Hyv9N�2�m�� ��D��P���F�z��xz��/�	����1Im�:�U�@Q Jo0��F*�f��/�AN�|%�$r�]1^7Br�u~i���d�8��p�]�d�đ��8���m�ɊMm�h ܥF�,����:'b�Ws�>� �E�GH ٪����93��xB�~aw��u���+K�h�+�'T2����ϊ%k�����]�Ў��?7�	���1 J�	B��I9�
e����wI� b����ϲpYt�։}�ՙ	�^zQ�� �;{aJ>L>�'�qð���t��O%6,>�9
��X�t���,�=�qF��
6/��fU��<���nN ��i愁�ȉD;� �_ٵE�3`D'�@fQ)ο��2;��lj��������M�d+�x��ryh������δ��d�7g:Xܥ?�	L�W�P�/�}��{ �U�{�|j���m����^9ͷ�'�+h1R\�s��Vs�#�����r�����!��z�Ɔ���ƮY9}���P|���[}�3Ŕ�A����!�'|b:�C"O���'��5p�r��S|,�G�V����d���,^U��FwC�B:�.ڍu��)�¶�<�x&
����?i-��Mg��ص�#}�g&k'����D	���'��#1�L`�{̝�`�|4ϭ���a��,�˫���B/��g]������lX�i	n4��Ul�w��L�"�v���-�y���]�`�Ϙ��3�8g~C<�')++z�1�x�)���Ώj�R�i�4��U=�k�g: ����0���B,�_ڮ������\�T4泥l���T�B���A�)�d��"*��%O���kP�/^�btS�U�)�Ͽ�������F����h*�D $u`�����c���xW��ƴlL0��h�a)
�s��;�;ä��"2�טS�2[���aX�y3� s����x`Nn���S:���rAPsY3�t)��Y��7�څ>�w�RI����@qםк�ک��_�%�u�i���yd�������'�S9�hgm#o-MI7A�k9#�9����~��Y��YcɘO�v�pza'><�5=R��B��k��}�>�J�R�RA�f�B%���>luR������D��m4������l'�K�Jء���9mY*�&�9��ie!ʎ{҈KY�z[�t ���qh�硄�*NM�_}//����3�.�2�֋5�'��`#^Ly�~U|��M1��S��i�����ca��ϩ�S�>��u�#;��>�6�ry_�y�#G�(�U�@���&����2���c�Κhymf����[b���c�K-m���_���$+0�����RPk�ʯ����Od����G�q'@�0E�`���M�<�`�_��y]|ܻD'��
8Ϊn�� �A��b<�MX"(9]b�shdl�Z_2�xZ*U(�G�w�ai��3�F���C�C(Wy]���-�u�"��t�������*�Dw��Ʉ{��<]��r����sh�w�p�����15�u�E��e:��]���r�I�ȭD&����xl���ܸ��L���_B�ȯ'(�k�z�R�]#T48���jx�bkg���w���^hݜ�����vX%�}���ߥXcG0:�.�r��h�4���4���l�O.��_�1K���kL$�	��~���If�
Ι���;N�v8b��]��J�v�X���ly6�,�a�'$����,�����s�%Of��Ef~�"�s��h���X� �J�C��I�]�S<�V�c�M��G�����K�\��mUwoi�l�f͵@���5|0J��uĚ*�v��צ���g^fx��	)��?���퇮��N޽�m]o�CYw&��Pe5\Ep��f��\~y�+�B�\�!`��Jx��]
=��f�VÚ�&��z�ֹ��l��$^�M���q�$o�mOj��B�-P=#�X�^�:p~R�V��d�G�j�+��gko׋A��k$���r:�yRr%0`Ś�Z���Ed��4�eX�]pl�|W��"���
G�J��j��M>6)�`C?�~ �5o�O��N��	�V�۴���}ę3���ḿW�i~	kV��U�B�Rad2ِ>e�J�*�h�m����~)m骋Wg���]�%�]SXX��ˁ .��b�.��c��:[�/B���D˪K�E-���qS:ք��j�������z�����x�8��ĸ���Rx���
@��	ggԠd#��t#���3eg2;�8�"�`���Y�i�a�4�&�2������ց�Q�gg�G+�6�Ҳ�r	ӵ����o⇓b�}�^"�$�a�o'�81.x��Lb�ߢﾃ�1i�%���d�Q�B�pC*���,c���۪�p.<Y�E�p�TU��'���퀧ԛg8E�(C���X�j�>bc�q�2��C�Z$�8h����/i��א�� ��z��7����wl�|��5�.��F2�\4(�쵟�=U�!�	���e{�e=U����!�D��t�|��}2�~�6�3|��2rZ��! ��ޠ�,i^VK�o�6ݚxT�p�;�ܜ��2  g!Zً�=K�pd�_�kF{%��r.��я?�"	|��+�P���I{�6��=�����ӏ�ۿT0(U���wfG�ԜV�Z<oG����;bqx�҈�����[�����Y�=Be�OX�^B��sٲX��qr�����*�� aK�H���{�h�{ ���a�/�Z��۰��t���	d򈹫�x5�s�!��v��((�B�2# ��'z�W�b�|�nyQ574u�?��>�aA�u���gL�l��[bm��o+��GG�K( ����$Qj>s���>�W,[Q���#\G!AJu��.Cѩi.M	����i~X�K���)��f,l�����]Te��:�p{u~}�XXp��殯 e��Z#�0��[�Lû1��<��u��7�'ў��Μ����MK]J�QdG*"\�U����P:��?�iž�:J�q�Q
'&�[�$�VQ�G=�[K�2�I�Df�J^%`�>姼�&�R��>� ��d&�wH�Gf7����~q���௑�ve��i,�[�r]�.ګ�Y`��������q��F]g��]��^���
���B*�˒"�BW�x;;�y��\<�_��D����Å�R���Ui[oח��NA��I9�Q-A�\��=vF��-�����¿��H���6�C�<�rVA璎�ҿC1�.��T\@l�;�J�ϊ$�:��ȊU��YR�vb��%�!�X�՟5�ZTR貔C̼�K����d[F�=I�u�N�ok��<�3�E˻����J�o�f�5��Ao��.�/#KN�f8?�r�ؔ47A̧�*J�k�E�Uݓ��w����'6D�OPg����V�N��r�tؐ�%�A�=oo"ӏě�0흛HB�W������`�U���~�y;C���\,���Ĭ�܂bte����.܁Z�&�OG�����@����w%9�ϒvwIU�"��ᴤ��
͈��ۘ�O"e����G	�8���sjJ�j�\Y�����ݧr�HS�Cq��;�A������,� Թg��.�$����4����G�K�%l��YTڢ�*�;�Z�fZ����!C%o�Ghb�Tja`_$P��YH����C�zCp�(�RR̟P]փ��d�.��<���|�M�'�G���h�(�T7�Q�9ֲ�ڝ�ٺ�q��1cI[�"�݀�Z�� 19�X���Bs�6�Ɍ�z|���3�Qm��m�ƇT�o�c:�Bp�M@�K��c��z�H^7�C�Ap��E��,8�nQ��2/F)��pC(���DĀ�Җ�V��  D����K�HRus;�J�� ��Y�¯9���`��XTm��? �5d
v����ߧ$h/ZF���ʎ�+�\�ᱝ�{3�_!L��C/=�Y&�q�+��b�o�S��b�D
��' lW TM�����r	����[�]g�g|¦ ���	�x���U�P;���'7�����(f��c�ݵ�R=j��E���9�քPo��6� ����fQY4�<5C�0��h�T��zm����G��O���%��N��s���h���ct�A^V�`֟2B�p��i�7yO"PP~�i���+@@H����(e1��ϙ����*?��>{L���"p���'�jT]Xhِ�Yw5�^9���:*�,`Ké����"MI�������M�9#cFֈ����P�L9ܸ��'N��g|��gv��3�g~�Ll�̲�	2�BEr O�"i�ɆQ۔��t��)� ��gN��?!f���/�G'@\&�\ǵ�om�u������ɛq���o$��
�1Ɵ��U�G?W$���sVc���&D+�Ht�,5�=tN�J�%xde�Lvؿ��¸��ɭ���v,���K��xLvpD��Z3�foF߄9�,��A��?%���"",��C5�+�8�TΧ���p�+y�~�u�Y2�Ū�z�Kn�0�����Bd�3���~�*��%���ݣfA�����-��E@G�z�$���,�ZiqJ}.����@��za��b���@q��*@�wy����E�ݒK������Ή�Oc��fA�d�?L�9��<���%,�g�[<G�����A�1Ų�B�0)v�����?{���Y��)�'<��`�>'
@���@��֝f�$�ր�I?d���b��8��wM��E�`"���~:��̑�`����U�M�F�Ns���Ίo���U-H�	D�]���d��#r֌li�A }�T����/K����xַ��W& H·���Oa�5|w6;�%����1��d6g�t���ltC�Cݕ1>/hRm�V����mbrv�����qr����
M��[R��ÀW�<����ϤO��>�)9W�5��W��M���M��f��_��0s��p�n���
��`������SL��k�ސ;1��x��&!�8���:��^��Dpo����N�Y��&B)yU�{�}PHAw@�%��K˗2h̕&>������1_pР��a��G�x�Qf�'J� ����O�\�5�A0 �\$�.�F#�R��8eC�ң�v�~p<��>��Y�ߥ�EŶ�{����Ip�]5P�K�����7:��b���Z^��Zܯ���:��x�)�D��Gdw�ǀ����N���r�C(P��#��)O��v���ʽ�9����Rs���m�3S�(Dp�r���_��{��:V�4u	=�j\6Bz윶�h�f��֛�a/8N]Y퉩�X��<��j򹋕��BPv�0���D�*~P4~���	���}���w�D�Ό���<���w
�`���I����|��q�X�
���}�nY���J��ۧ���X�4��Q��9"�O�@2��� �(�jp�R�~b�?}I�k�����~/req�C���ɳ�?�獭+f���mc���/Y~y�wՇ��ы��Y.�W����^[L%��Ԑ-h�y	L�?�jt�0޶���*�DQoz�A�k+'�լ=��\�F��O=!�#{W?獂	xZ�裂����@E�,���:�ߧI�p����t��}ԏe�aD��\,�J&���� i  
�b�t�%r��so�8�!�����z�?2���Y�s�Taá�1�ȣ��/d�uX)���kS��9�t)�̃@qU�A,���_B9����J�FZsge���c��sr�0Ұe�У��=u��v�T�����Î���`B?gU��.5�B�e&��x���λ�`��e�7�׸'E�W��¯'3M�R��nV��Lm�d���E;��T\���}���K5��`3����%1W�0�U$G,��墯h,A_8���	��$B��W򩶦�����HoA������Di�G�{���+�=�ef5���d%Ͻ�;Ȼ�4r�����V�>�O�EgU*ܳ�}$.����M<����EXD^�r�� �~��IP;F{��v2^@�2���赌�~���*�ИؤR��$��H���%�"�80�5���g�����Tr��>�Z�jZ�u�~�"����]L ��0��^��Z�ߙ%.<��Ko��t�9�;�\����#G��FGEQ��c��f�����"�Cѡ�*�J��_e+G�l�'�Cl@���by`S<�aՕr-=�nI��f�@�Z�B{E��u�9I�U��v�1MS�7���yB���O����33ݛH��q�H�=�2b߉���2(eA�T�}Fr���Y5��F��!��M�r�#�o[E����qX[fM�;���o�ި�C��@a�E�\;��p�\��$H�����OT�9N5.����\�LA.���=4�ֻlz�%U�+�c=���0S��le��o�k��P+U�0[�h�d_4遽Y��"��«8������J������:��S�V�ŋ��*)V���T��I:P��M��[�:N}�oP��᥂`�x{	���s�\Mt��8V*?0c�'9�+���G���> 4a�L�џ\�_��2l8,���`�j��2��XY�y�Z��F,l�EX���H�#W0��B�-=M�5zj��LNh2�}k���yƏݜ�N{��uC� �-�~���Y�H����M�l�﷥�.K��&����\)�43l��?��H���	i[�i��(��G�J��
34�o��:�aԚn����g�ׁ��)~�@) ��`bkxT��</p�Dlv �J'�� ��A�r?�,�!��|0ww�oЛ�'Χn��� ��R�$�A�U
��f�g�?#j��	"�]-����'S�X<ˎIӴ�[�vk��ݐ ��2�iffk9c�l-����Tfb6*Bpo�^���)�h��v����8)X=��:�V��e����GZ('�1�)��k�?5%6���l�<���Y�*�a�n{�z�j��B鼄��c����;���ChN�P��~�.�D9o,���T�+����!����:p�=��p����?����z#B��\k�{w�Wը& %hs��t�B����'��4X8#a�{�.w>����Gʗut��:�!k՛i�9�>OiK�7�i�$ðO�t�5�;mW��`7jiG�bc2W��s-]9޿wz�St�#'��B, �����d$e}RZ`୹��r�u�e�����H����[�A�a�8��=�j��]��B�u�H���CI����v��*]ca����ql�Ĥ8ۃ�y�ᨹ�So�v@m�U��k�*�[�v��~�Hde���U����g����M���tj+=h�<����*�2T�<���nA.O�ڳ/f��ʝu���-���ݞ&|�$ʾ���Y�t�'	&T�UΠ���q�_J�]�"���)�8�0�&r����Bc��