-- (C) 2001-2016 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
GSFQ/xXPKUwaA9nLDkID7Nb1AWF20DUYj0kLQ8haufNub228ujS9KE/IcCjKl5pD5n2HXpATfkmn
16qZ1+OR3eAY5yLbMv0f+0dNbvmfnGbGgu0vHM9qgr1thWnU3Q8SlwJWTQxOpiZq/qrjsdT6ieW8
VvcsCiZT4Gi45UpXcHzRb8vwBfon7seFeWhDEAHj+BBlHVyipIFB76a8udZnN9VXPkJAzMxzEgSh
M+5zYjMDGfmOf+4cFDRVQXfuuiyPRZv346BmpXRKp+XIBU2nriFuGmtKLKDTIriI0pbgxqF/cJrA
mHbg8NruYtl2/KjaQDT3XCZ6Cn0fE4UWj00D1g==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 6368)
`protect data_block
srHYCFD1nLl7Le9vZfuTW5/u/2XySdZ+EwcrFkbJnCV6+PofBTKhRbKikQ926ZO6Te3qN6gis6DN
fdnnHSRsgp7j2LpFYJ6MxXArq1hqQjJDYg9e7Ubot2sdJTxLBs7Y+t/2ZWb/EXqAXErPodPm7xOD
nI/NI0dmQ7xPKjLnkCZ+2ihXpLlss4XqLTtOstY2q7o1oH6z2dPucmBJsM2/Vw7ra6gAs8X/Vz2u
VHniZFI9/6lR4Z0T/ammumJipsBiBfOP22tHaxhKbqXud0ItQqN2/4nYAvHFBKqn9nYQQp9fDBPC
BIFw97TR9LPy6rnjjiBe/2Rh1rBthbpNGXESpE43xwIMib9Gdyg5jWKV3/dbCr13fugA49mWsZ58
cBCtN0Mc/0ZAzYJT6fw1TNeemDqcQW0slBbxJtqzdW9HM99GOjB6xxzkosZVIrt1K8qyLb2fzxXN
Zmk4Cnod69yWBE+MhjJy/Jty0l3csb9tJv96ipebrMzbI4qqh4NsBBDmUXJzKRQVqqzLqkqB5SBv
M1oqP5XrFTSRysfw08qaD9JDIOMqtp9bTxjKsQedTEg94xuI/rcBTuog7blfjXTZDf+UuqURaoig
Va3W9pDtldQJ0KKxI/Ny56S9jFghtbwrvRXqwsEw65+tydVfXJBg6LF4+oHma5ku3/vA8Jf5tvwM
0gGpklhC2dS6rGUOeCNti0fSB46nz9xAAqfJaUuQMycYopbmYhLb2LBr6ksl/TRzOS4dmMSbWOw1
gi3yjxcBBM29v98vC64xdvBR27Rm1ncxv3iDxOkWxu3l9JSjBez5NjE49+EpPICIY1pxQRIU4xv3
VM+ATU2DD5bRAFPTWe/EXgbauxkoGyfNWE0iO4PCP2zvYxX6SlwNowNnR1FHb0h16ExOodSbnbDB
bCD5eoAsiVoVVJAQRv97BjnjPoVb9/cczrYHugBsTSMwgo/exZrdDJOAnZ9e8kd9PjmqeRADNwMk
Wg/UdvwwmiChqSJEGUIBLuzmJ9fMWW3lAJfsVn/UONWhy2VP2rABJZmHG3LjrqvZSuQ9nrkrVNDp
D27w885iAmsx4/kJthyOgH/0TYi4cNDcnrSvqvBl1asgaWmRrqYNbKsBBm6VyRX23Q8F83x73hHe
8bzFJHXs8V04zB82mYJ3DXNOyFiHog3vlkMZscyVb7fOtj3xAnWc5wTmYbFJkMZDVs1IAmgGiDi8
RBc8Lqx2qEKavsdhrwdlyw03V1B5LtgANwSZBzK/ruOmbYFS8do+PkFwUzuTWHCj3SpmhCo97VGH
xCV26LzqQvrz2JHPjH1MB6mhGEjd/Far30l+8MQFJHE6TfaqTj61fBtbJ96DBQDMHOYzDZ9FgzHu
IJJ/mQTH+vrczgsZ384PkeocegHAWcxDOta4CN5Oc8FAr/DLPLpcQ/dUPLc8c+R9VIV2OZst6lHJ
KD6htaeJ1BXX2eFY1chjPVGZBnSF1uHEmpi15+m/cVphwxf1wKtyD03M06sN2/miy0JGcvP4gbtO
qXgkwYCHRWUVn8qqg4iUikj6GHKlQQ/DbnMM84QNTL70cfgG8OqHFj9eLjs5/qlMqUTUr0Pi5+hh
g2VQPo8uhW3YRKLVT8yHOMSYkG1e0c3anLJEzeMPoasEsbO84zHguQf58K9wf2bZ31Y3nFE1jG41
l9oOpmUVe5QePepHJL9dmotu52sykMLzGlX5859HkthNspx9WykGTOQopBN/JRlwOBHYxz4mATH4
owzNPJ7hGLsTti+Jv8MssY77UFVyoRPs8NEJ5plkx/p98kCkoWiMcvZkSXqmGpM73j7fsWyvhHkR
R6lxAOo1rzBNLgSHQp2mopms7hmnSXyIAnwkoDiFNYvhFAH2zsywwC8qvPrmWeFyInBg02VeANrW
pUyC7VQMMf13uiHj5mQKgsshHsQ4I4qX+/6yM3sOHi5MYFvFAirfZHPoxxX9emOPFZOBARBFEouq
oWz1L4D5/U3QWQvXmc6J0Odi8laCfQQlMvyBDG0tBPC0vbkp9JLfJipbSs3esMv9AdWlwpFYEIfq
DodxTVsER0bcnxPz9QBvJnoNDeEIuiskptjslcF/5lCaM9tmECK51DxstCDQ90z5C+9VHXXqqCF8
rwSU5qjtHvllFKrei+RymyRlo9fSK4480ybLJFywSwJplS1vvE/OQhIrhl8MDrgEOwo0a79U6iG+
Gpnd8GDrcIxjq64dDWK0IIZWAtpsH5jEAwlzWECkIbzQtVEIKaAoiIXBhvEnB37tFZCPUMqQgRKy
grVjDCvW0/tnn6sOCaLWvclwxalpGf7VW6OzrXesUkjL8sMJf/Z4yyT8U0L/dT8i97COkcaQBHGH
P3dbVsUfwWfhdsuVUKwXTXtyCBow9ZX3p45nJ8yTwq82R/r78kwcGnAmOuhziT54E0PODc5ZwEEd
8s6fk9HJ/Bxb+8lF1Jn0AJOCLXeQdbbSe89ky7jYDBkWr+nhhVHBIsuKMO49ZqsYv3cMNDXW3sUH
HOi8Q587IGMR+Xk0fgHko92HFknaPiGdSyrZP0puwGCuQaP7yAiDahBPB4Muo1Q+dR6iaYexUDQg
CLwwLERcXISUtvdg2nX5DrGHJOO49TFuvUNhawaYuTmQvXI94XQu+x1bC0vOXMjdf3jrrstz+MMB
y2nsIn881Y4+Gl+9dN4QDgcw17qrUH4wgoZvFcOVDQAoAZ+DmqSJJkWnPEKq2+o1Xqy/ETFB//ZF
qEXw/4fmmUUFVRc9V/pcNKXcYwJnXqaxE7N0ftLX53auePHhm6jPeKoKF2bF207XFwcMHBqB9qcV
sJAUQ15YyRK4W8y1KQHEl2f9vP4guryNP7a/UzhlA2PRqtJgTJYONptK/2acF7pBVvgoVr+at0Dx
DXhIn7E2e/1QXuWv5+XT9OJYbJVF5IOu0J9iH4OQygYU3DRB7D/3efYn+SN/K7LgXzTQQ6e6yyCb
MXuhKHlN9V++Ik0/tRpj8n+YDO6ET7wzPPhfQ4fN669B5vQMSq8mW6h7pWcydW6SvnFe9B6aK7lc
WnbMgKhVf94Vd9UdJx1A3H7CxMWi7s/13PUbiSXSSIQ8ft7Qi54eu/HEahdjXY7LqORfu6HsPt2L
Qd9aAEXu0tX2zL9sVqGqS7JpgTFZMysoNhfEIvbkbXhFkihQxtjZuX9M39K0W00QyocZzL6qFhrI
wYrm0b+ZhjbEANuH8YLWilC5/QYkTQA3Y9IGlXs0kS3E+88RxmzQApqx1LbVn3sBx9e+vOlFq6Yc
WflgcLbqqpyxs+vLUZk47qFT7Seje9O1TBeibdDOVs0B2Ba/pdYWGtDqHHwrp99d665NHR4/ZPYr
G63KWQsbybWnUF38tTCkzEuh+i/cjnffcPPanFiLJG4gh8nC1s3qMpNk59CIcY8hvV6EVXYJbxpv
y+N/89jSMCdZKn4sZY+dOaeQAh1pvEro7wy+708cujl6eFLisUPFm/iRXQ4epSXgkXWTE6zHWsAk
Mr0x35Z0LyK+wojFXqrQNjSyhw59qZchIydRBdL72CFvXsSLOAiVuQFtc9VQxDjgMxqbdO9UieeZ
89pgKxIGaPnun5xJghpPl/PART31k8BFw349wghZpgUQ6XlKEAnkWSMjr4w2HNNi6aRR9lkRyv7r
/GPsKmunzTjjFK/HckdcM4pgquoLXEkq3alN0n244qfhnoKWI7xJuhTGHoeEkqn26RhZHFv3iN8Z
7lTk5XvA0BJSYQtotDuIihsfkNlSfCAqBxmHg42hssCHoHXuVaRDmeCkUlDKxskvql6VF9yi0DS+
8zDmpjDp8kOBlDORY37NUn886FX4AZF+AlzTfHeJq31MmT++0vq8BZ7G4B4TqHNmSHkV+M249tyx
M2U5knIMB4L2ttc6Ow1ZBEdqD/ICbMclD7IxAygDtss8IRdr8uQ/Z+SxFkPNMAV0QN6I2KcvU6S6
AOg4Vd8qIIk96G0qRJdEcghzj0O6vS23/AP9MRjOhl5RtmU2vM/qkk5iASTD4dporA2xJuu093BA
gxRTX1yIgArNowT/xsd2m/JeBu9Ne+R11hRl5Drl4zDHf0/uwBJ5Ghw3CGvOOTEPpLLor4DO/uHD
zZEiv86dd7DfLNWs01hhfAEbhm4lMz0/yr9DqrTWmEmcZxgu2uGOV81phJ9GbQU6OPOIjr3nkjpE
IF2jI46otxtRYpQ6/mvGtw9zJyiZ6r1gPwtMQR2KIg3gqlpVpEiQZkUZKIIqBdNqJMCFeW1eGEH5
VK5wDqOdk4veL/tlb5DZoEdgWQv61CjfTt2mRez9v0ktd7u5cNw0LLw/WvM3a4WY5u1jtzH9pvYH
7baGVD1yTymZ5+RpslKQlT3aCZS/VmUrEwpa6X1G97q7nqYOyt2DAufSidHuAQYUEvB7B0NBczuL
1jrZuk9XuulXVAVTAq4sqG7PbXblFuVo4AR/5iAdH6l8MTmv71grols5ePKgu/sktr3g1M1QRuGq
ZENGXF+D4g7/UNq/UxEE4YQxAyADfOFJBsHBHBBT2iqlunyjDHBOBvgHE6cE21p+rNmsLqo2wOz2
iL18wCzPMDL5D6fQgDNzRpJffgFwi1g0wBmTO7wapiNUYP6oGI7PYWr0KpIWm2IXqA13+D26XSL9
TdaRpn4RpV0G5jKk4VJQiMPv4d+sRyCT0AwEF4bbZRytwrroX1018UeuVDIGYWV4jJiS5XcNr+13
ar1qYn3Wc3JxKS6b1QP6XhCdkhi6EgnqsPZBi/Y/NHTjDs9U1xfzPYemKSA/tfhQECyjZUv3IFdU
sW/jxI0DDc6i2KTxMo34Qkjov/s/YvVX67N7VauRod7PmjoXZkrRL9C0FjjjY/jTBJyaM6rSYw+M
kiEZ72QCfgtscdL1mZBaDM8v1tWtezj1Tuwqr5hfZByJr7WGnjdTSZ4U6pbaKxGWbiXZzHbMO1Yd
ldnJ1979pVIXyxnypOBIz0Pq2szEzS+xUt2ldhxdgoY2G3XOZrbBqw+Nsp8rtV6EUM136MW4jBYH
+y1nZih+zzXWqH91dNIKAsnOyGIL7suJ86mVyHq4LF6Eedfa/9j46ZGOvREjm6GVRT2Y/7vhfvxf
1CvZe3l6u+guDaDE0nlcfP+H11lO36EE4YF05tPhCx3fc0czomeSoMGqs9J4gx/bZOxu8d0NPo2q
MPqht7ArNm9/F6sAj9iZzsSjn27013Zg+KWQDU5lhV83Ah3ZxUrVW1ZI59jx75fQMcKCjN1Gtnb+
U94Azvw+zqhvBlXjM0KO1oZWFkV5YcBGIhFTmCwesVIHghfLsqJnjz+Pq7WiXJOGTjlKkI1mV8Yf
5VP43cKNKPPMvx6vCHnzjxClmmjfdKWqSFlrIWS/EOYYF2bcv84IRvca8CUe+KN+0fF5lXCQYUAY
jWAXRZASjUJj7rHOgazSqX6CMfL/dETojtpScf7zfHl3Jquz5lzSdx77iyf1BgitpQnrFlkXUZQ/
GL5X2wLZFEDcsdGbz7DTdzEhUBpPYM3ufFCXeqPqN6IPeZbju+nnKH25JTHzeIQAfuPauvCMc3oa
7ANvmePvl9Vd5eCFgcLq+SEFRqfNzRaNXODAZgb34lPsu1EFO0i+vV28CUfkwq4PK1Siu/Bd7QTJ
GlMeHm84k2+feyZo79q/LzMACtF8fyLMIf7wQLjNPdFuQp/CV8sEweafibNZlRv6gaJyJmetj/DM
NatmKwZGry8fK8VJR6CaiktIefZq2vXLbHvxHwNNSfp7DAFlufJttdSNQnEXeRYhrM20H341pNrz
ZI27ol/nRNhemEDFWMij3v3kXIVZyZQ7lCjw06biOGKuj4o4Xgv8zKN9wwhSpDfpWjiqFtaNlzYy
6WrTV7yjPdxXMgGbPSu5rESau+kfpCAGonSDv/LVaB3Jxw4zm+jRCD8HRr/pwZIyPqWnrKzKkFix
75Yxpzs5+qcidnU9icNogga1PE1Xeu2rhb3+6F+EP0+cZuUTkN0vLG2iVwpasAAzFN7UoXn626nl
C5WsCPJNcsknH+10+gMuWpzoAdjG9+8033jVuB0Z6C/8ujATqTdtpnY/k3d56PWC7+e/KQ7PbQEp
0ZLhNBqiV0o6KYRa+xVShTcdeTF0g7y97oiHubJ6GIqIE+cbuXGqC65wXcUA3uy+cZMyqy7zpUO+
DcPuXbIcNqFBKQd8ahhO5ngMOgTfC7VesNWSCyQAlEML5r2JNMbjhP4niwYo/si/6gsEmLlEXqqT
wyL7nIrL6apKy+EWSw8YIU2ntJpMimAbddXgjeRODgZViByNsikxHeUIL5NqeRe7fin8o4qEWLuz
iedToJ/CVCDX16puSv06VY6RDTAANn/hFyNhUXIYYHOzxYAruwVwEmVUpVJbcrIXGoA/lq2kKBfl
QcUmNatWo7kthckXgS/UODasSGbN1w177Bq/HD1p0ZSbRY88Xokltmvfted81bO92gCdY04hf38e
QyiioIauydo71TDw2vqUm+26UhnKAI3Jih/ZlWX2rseljcEH6mZTF00OR4Sq03rrq+lNTtbVLfgO
qSgSrinHDNsRpKQwlUUlMA5F/EnpAt+D2m/f1KNVyRE0l8yQywKX10K+ZQRzyseuIEpJ+uwZkL9U
YXUg3peSlqbGU4d+SRML+9F9jo6f41ZCM6OQdASV8BePHsiIwK5r1MH24NWgr8bncfNUTW0coILQ
q2z7rpRXwohdQVI2NX+xx98da+N9dEolvsE4ztFFeangIeK1TwVtt4xVJl0ET53QIKdfkXoVDvhe
CeL7Fiw0ghnyDM5valnUCUK39PF6OlnVwiBaSye6YOhxLL+IT1fvlMH97ic3oTUyHV1tTB4H2VUe
HSn29tmDdlmAMofsTEms1Zfyh2DZXtivJrot4MNFzCYB7rbU+GHOByK89j3IqglQWxLACsy46jPv
TzFnZGsK99VTbB3AubENhEXUc7toD04AnzHwwNO+QfDPPWBEGEEYKuosFobed6rX83TMyzjD/Sml
HnDxtL6DUQ47V/QH+4tAHrpakIlyEtVt73rdOUkxql5A2Ju3nYFo6fDFDbJKK9iykfoQbTeTCvB0
hN4gjneNuRaCxbf3cff1dmVGcTQ4BK0R1v85W/xJzvZAjWuMciwHEgwvrJA2/hyYLfnjHbFL4+eS
1cI2V7Xv5nXOhInT/gLk4Ymnwo67xZ+fM5s4VA2mJoB1HJJ3jkKJElLqV2GD9dzWGHVYEo2Ni6wU
mfur22jCSCzT9c+t2mg3RmhHNzWyhK9gk1jOLf2T/GKIL8sm5b/oC2Ofz5JTPAzBEkurfeUL1eXi
yb6eJTCUq+KVLS47xJArox0AeZ1mrZj0PjmkQp3Wp79iMY47zUc1Tr6GzuZ+Z0VAWZgG67i+FSx4
VfGef3R7lqywYimiD39ZV6qnA2as7LxN6nwG4mvCKvPqlwnx9Yt2E8l/SawLaGGMTXEo6y97Nh/s
vnCmguUTvb0r6uroM3lTZ2LwRhCV51gkpafaf4ycZ+y7iwbqWX1y1BsXOPiYjbdB4J8lYqBnnLfh
0t+Ua6Snzywgzjuqxvh3a9wARrbXcO1QFgHjKUFFfpevNI5CDQmHXx38Zbn6Po9X5+A3QH/eeMjd
2g8hvykmQj6K2R/qOaQTManeys6pGAmAy6uThtG93wBsiICMhEQkoKr1l0OM7w7J7I0c/BZVrUFK
IUlC6RFVz7AqV3TrsQI9UuZrEuMkqSDu4O7zT6e4jiDWsTHXZ1bZKJih4xNjNAB/vd2IeJaLs9gS
vLgevPi7tAZAduZfVL3ClqbdELbbtJkFN/BA+AjTuSK1eDbT2euvxM8WnmqFKH6IVLjDngjf8Y90
JUEJ0S1cl9KK+C6oYj1Y03xvIzeWGIpRgyg8CGh8O96a3MZZBxXKBCbNWH6359GnmFK/2ENUqIle
xZGbDlyrqMTTCVDGoYh02K/g9xP3KTjkvJInjWsmCXAin2+/tW3RD6BzQpbuvnYP2+IreaFcq9sQ
/KWDkWARExPaPG6izY3ftGQy6YxiexcKkQD07IXCafvo7Dz9Yj9FXWXR8TF7X8846Mjezdc7xVbl
pul8gbZ+6yX9DwQrZeMWeQmiigUdiQWGSzKWqm2Yi6aruIypPRei1uyNGaZHLMqjGpz8KNnkOlQ3
RmTbGJ9NWUgc4/bH19GoVztjZsofJQSLXSKQ34FnYJDc85YTCmgMDu+LzIukkz372vTx4Hfa31iz
X3HRkv9KPgu0hmtFajaruRn9mAVc2Gccey8ZawYkJjYPIPCdUJL6Wby+OmUAWGB3vrjgvgFhEQNm
o4ORxaHnUJdxU90hco7vKyY1TJWcKNVtWm5BM5GhZTTh5wwRsn8YES3Qqb5p60KiDSIVckk9VeV0
e7LSN/3hkIJ1Smc9VWgge0mZgtzNlK0sU9HPv4J8uBfO0Igaszsgmy7eYyAyxaXktQX5tK5TfiQ5
3C1jc5YeAfF63GTab50xUejep5WQ203QxxTSF0Z8rEmhTg1QR0gk05k=
`protect end_protected
