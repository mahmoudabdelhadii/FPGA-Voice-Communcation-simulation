-- (C) 2001-2016 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
dVNz2iiaH7yvW8PGQNiEXaS8T/JKFMLhDM6zEjPuyAqRDN3iSUJBx9nginhFOXOL3Taq5ajwjN2+
02bAMAuNM5bnYHaMIcKWYiin07vsLzgCin+wLgiKijzrx33qeApIDVdOietWxeaaxIY6EBwO59TT
8bNuhjxqRbThdMj7v/Nn9LI+RA/d3DOLbNcvZSn1UzUVHta+G6U+97L8dBu1aSvX67Pr997pN7E3
FobQQ75ahaEkF0IHTObX/iwJH9Wmzo3lYtInieHhtvxQ3c672XV+fY/fQXWIY3A8gnQ3CpFlw78I
JS9oczCbfDXH3vHOmqokLjUIc0MXAJKylXcgyQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 13168)
`protect data_block
QXRWay8KTtyj1QtkYdJGXKDtJR7WzOtH2qMJ29um/t+xswQF10orgwxCvX7UuIJ7rN9NU375zWv9
nRmIsFsxOaxUxVCRlxOKbiA6MZ2tLCy5Af4RmzU3dQ9UFTiVuu2lPtz3YmTzHgU2ILAHvqPAD1Uj
iLm5YW6Iho7Vv8qu9QsTFH9wYBt0nRnARi9qW9EdiMDmSrCTrQqnnx80dPfkGXz1+ob/3BD4RAiK
yokkgXet7sGCF3mro5ureLuVu869Pvr7mHwn7yf5x7DwBbgEYSyRIHuj8+E0chuSXZWphGyEBWIH
H2p1XLxPLWzY9EpEp8YYSoOOeFGPixheNMuhCZokD1RWdChftKPGqKpUiQ9Z4MvCiwzHA9oC7ugU
/8bsI1p22N0jdm9lFC3gv1d5lFqwPLJSlUwgp7Ik6RJdIAQbot5g3vJoIfA7mKBdYWe9SsD8L4SM
ZjbPPl1acYY8DAOwdlTvknRHjZrVXdHpQXieh2Sf5aojUQlEvEeKUQGFeUTopSW2g3akkJmlPWfi
h0J+FcEl2W4IvVNbu+RbJiAU/Da5axDnqrfm1Y6olkH8KnB7XHz4VUIB+b/Ok7aJR43J79eDgD84
NOAOccKcv7VB+1F0s03VL2Yr5svy+lNCAJrEvWKYWF7i4ZUTstKDwnmjyOTpeoQH+a1pnUdgpNwZ
Ie44Ezh3wQNX1JpXDQDk+lX2U9DIvlmSNeKUB6xIqN8gVRu2ZWGvFRh+XGvY73wNF5HfFOaSlxUV
MbikETk65Ydminy/4j3YEfJD/6NrpNAPg+iEOpXHoZeRyeYQx5rJ07vtuWOfNE64W5T6vOXjT6a4
mGnGuag0r/3FIeqq1N+NKOIo7HDT5RQpRZl1ZfuIMf8AmnXqEl8XJ5TsEcyNYDaSCs2RRVh4NIVh
r79hZKDjiFp4kVGbkbfTGjJt2lT/IdsXnqyl5/CX1l1OccdwlPMHpEAv0CVncrgM8Ku8efkPkl4w
hBb1NB2fEZmS/+/ddMqSpKpVTqASPSrf326+xch7wl8bkGWJ+B43FANNEYfqXfRZ8gxQsRDFqJT5
Wetq88qbH4YdnQ/UL00NBO2lbqJn2qf5fR3ebfXlMtCnj/Xov3zA4kCRlJrZY4Djf7ic6PTYKDHJ
9Dd3tPtF9IRAR/QjALOzRfpi50hUpNj/yncZIjSTeVE3PlSZ8mFipWRNOzYe5W6TjUc4TYdUnYyR
iAjcRc4F/SRN1HIeZaVhZCB840s/EwJaBUqtceNK92hlfGgRFK9ZSYZBJzMWwAHCI1WjHgpaBVqL
LBJGyQpW/B2ntgdSqQ+F4yUYD4oMIkT+qqMXcS5iiCzs6FmJYZhsXc8O/ZN0nrAQxbWcTg7RQjHL
ed/Jxcc3WJGowurfxL7QgAg7DUTyondg3RTDq4lQTA68dwkISTvHb2Iw7GhTJ6mBJriGa+MjStQY
tPB0yVkYj9kTEacZtNewcWMZF75eRkgIJwoaRbI4sr6CYnRpgLaqWm16D9b0TW+T6A/LpRdAQdk9
zmsjnkgL6hyOAQZDXlqJvLtSMyC1SWeAkzz6IJqC+a/3ImQkSegcX3Smo/ITZw7MrTcj1HdIqih6
dpOyoHQSNHCXvOKDPkmkbSkVrMndmof67ciGQqLyeTv4XH41SzM6IlmuMA38aidOAmPNsa4hSIGs
gsazkISWLBInjNPPsO+AZAzat3YszlY5oJc7vVDtuifTyEfkJFo//MK/fGfUbpe56iRTDWoedWpT
pPy5B184UT8taCyY69cj6pBuwzh58Af5X/xwLM9O+TsIgxSyPIdPvb5bDqaNsQFNSfcJNzyXtk5Z
evndqMxTNPIpdaeB2DGthVY2KFm0JGPbKDLJj2oFtEekJJXKLJq3vA555M4sDNEpAlqbZ/nNFw1W
Nv3prJ8IzFLTlBRh+mYbmUR9XZiaS7epLNkLzPE/QlSoPsoKKJFZzYlj5WXSn9RNaytfPeB32bGT
rFesxrzvQcCuN1kEuEzLkmah+Fsv8FtJ6nPkoZ+eLwp/yaw+VyiYBbIbZbOaQhPYDgM034dRfMT8
vFv33nKZ9yAKmm4x/A7Sh1itkA1qeG6KK3sQy3nph07W4xEdxILOTs3E5Hz7jbsi9cGzNfRcc1r6
/PvDSh3qJ4kdMLrapQgIAu6UGHuxe0fhTpe5WY4HiAj3J/8uiji0rt8dIhPHKwRS7fu35ZfbEtyg
ou6OYkGtTScnNaI8jdHNhmXSgt85lUmKao+o8VXzkLyrS09GAKkA+F8hyNCSScomTz9yGCGW7p/Q
TcvVfWYrAU9Y7udnalgEjL0qoFhklBgy3re6ouqNnB16qH/i26to+lHznyj4HfO8kiw+J8KNY7kQ
e0gr5HyiLVU8TowFN9NxZuSf+Y2LZVfxvmmXC/6fqixnhi3/94yQgsiEzdnZ2hREncMRzAy2aa7e
3WvHk1bnp3V6NlmsQ9LAfCXf9LoAIWvapVKgYHw18cK1vHqLsXx6Ghb7PFixs3EY+auf+1E7XLAf
//Hfqs2QPRUe7fWph4AiDBOVHkpuag0TWQNFtg7peX2Q5YYFypDEZhAfN2Ej/Ds7xGIPt0P2DZOf
w6Z/ln+L8D0u3F5hBxIfZ4lY8ot8EJ6u3KYIuMH5EEW1xBsp9GqSbGbmN7Xgra8ajwqA2ufS4GNi
uMa+bHzVjugjdCIa/FFY0U43Fi8l0IEKsT93Tb20LK4zmNakA/dHWJMcZD4Jq3LXtnPkPoYXLkJp
BqwQvAjoLWKZfWS4GBzJGp5NbIe21cjuTqjCcYniU6NOo5o/L2C+OQfuIUy1cWqR3Jj3eWyinNvj
jPiXCjL0V+lwnfoGeByFVa+8CmxKU1qCI0nTJIWXXEaiz8uDf5ZlLMF8HHwDjVLjAdNuT4N04kgE
zHgq3ueRqxAnjvk4ONeQNpdHn0RQqNlsELN3EUUp6JTswLmBqnvBytLEIWoG/ihnGYn8oVrTxNp/
1TZg6g5ZaBl5ho61Yj+dyymMK8QbIztaPFaPi2xYkLUBZRUaSI3MayB586RXTXWW/5OqfmLBP9kI
MOPSEUP1KdGDxCSl+iHJAR5XA7S0hQYCNrsa5PWPezGJLvUwA9c+ZcFwuzrdQ3jlhLtoXz0AMSz9
oFacdlYfxBsm5SwB0iwdaWYeZjjxjv6uTsl/OW2vdW+voXusEgzE1j6U7qzvzL9rkkbTTcJtM3dJ
M46VECh0jOIaStjHdrAjTqKCYMAegI9lFWEMDDNtm1NNYwGJsjFqTsdaJJZ/Aw0A0dZcu0+Cd/Fc
44eZzxbXHWrKYjJuIYsIOyBTL9W57VO6QwZwB9Hf/BrzCPNEwD8Jxv8bdNFmCwBXj23fdpp/MhUm
/HQJxa2GJeV4Lzk7fzEHAUxF8HxyJSWPrqq/d3skLsXZZTGI1oJR+NZ8vphjKAveAfIjzyjNmIGK
I3apaV/JTpOo1fE6KCC598gT7+Vg+8z3VOcrnOuRZ6adDUQYFDBxww5uy4MAt8tJX4gqgOF4txGs
X5WREaueP772ZU6qBLdqqvVsrO3jIqeVkyNJGZloB4xNGlvyGt3Vo2IlOh13dOaVNIgRyOognklz
iPbmx9ZguPIWldiZmUay1DmwLtbcXN3WjOHaPW92rwkvz0zYf2Fgag87T49zbbC7jM5HXObMLjws
RL7/dbpiK6j0bnVNWALz6cMsQG7/z/HiPYuHBZDpTABFmY9gQl9cCKgmj/Oo7vMaOpmKlvMRurF4
p4/IUJF0W80p3MRTmiRDaCfYvrLX9Zn7Dm4UH9BTK/ksIkJeOuMvIx5YRdZx0P6PVIkrinhFNAPD
dwJ7tqmofsUg6AoqLMKQ+wzhr8/ILsb0TMwqigd+7KMqSiLmb0rtX/fiFIUS7JLSt9nzPvKuS3Fn
AW+TqOwhwLAbhdWL9SCZOlzH7wwEJCw44535B7drViuHj74PDKhHw4N4dbM6KzGcWJT+oGvwKjDt
wYwutS7/E8ZhW0wOSc0c32kA3/EI/azlVguZftUiEzwgR2NHtJBGH0eEDYzX42Hh0FX2SxjozFlQ
FGKdt2yn4fqX1d9vFC/T8xd3AqDEd3BSk6CRooeswjfjC4Bm5ASUQ8Ej78G5S+JIsH3fVvct7liM
X0+r6HxGnMFP/C5GotnUlJGwJSo9Hx38JddJn4V6L245A9K4GK3xa1MEpRR2hOljI7ozpDGXu7kB
O3iR8DkhJEGKrxJRE30Y2SjUvZSHAtNoEKG9tK5iRlS51x5ckPNjTxpaw6KtMPxtbtZC5acne2Qd
8twUUd8AJR5P9aXLaDM477rUnvJXYbLH1uPJ+222LKmRcnlZ+F2S7gvCbtL76IjHa51wtU2YgiUP
E4xzEyTTiceDJKR0/pVpkMsZCdOcWmh2NbZ+kOJxgGmXsWtGVAIDZ+myZk89N1Q78+NTHdcf1b1r
EWQfX/JMZ2mT/DaSjOukDrib+JDN61WoLa5Fc042Cll0Lw9hjGPmU9faMgG45lXKq/KyrDgLCYoc
j62lNX0x/mXkiVs1oYMyxx5XDrMm9ilQGixSZNQEnVHo2w+uk8idDRuXd1oOLEbZbWv8RHpHehgK
FVVHADmxpZnPtpnCmvHnO+U2ajeKR1ImAqfwt99FbNITfEoFY1OUlqeQt2bwzgmgaehomTOTMEIK
XIogBTfSe3gjzbIzi62rTE/V95AV2EcCaNEf0rW3J+K3zvEQTeiiYv8bR44SoHJRofxXCWavDs+s
ts4V+o0q7E0r1zmAJXFdUf3f3wu2D5OS1UnRxspINed2Mp503IJUqhYCVlTDMjet6epOX6RUILWA
BcRWDSE5X4wRO0R2gopRtlRvPkn99JWHRor1YkeEzLQujcbK7zzU24umnGl1/yyOyUBkbswUlENA
mZSvLL/WyinKtTCrJtSq6jzkHNJ00kbsMRJ+ZQ149v5pJ+pVJpWFRrJmw5wpTxOFB3iLRH+XINEd
R3kVnG3XXv2PHBVEFLxfTcT6kd4vSNfv90ah32cFB6o0uz4cVyZgOSLJNIlTvJW7jqTHyAbhyLhh
ihN0oIaHhlI9c+ochUEvBgoUT/gGJGoZHCDW5JOuGAClrJJABwqeuyk/euQfPGUJNDljjGVMCjGP
Ksp+LXz36e+SrHoWXaXLpobVHSCxUUWMLEp6XDTugymOBJWkB48jnsuDEKm7tg3mONPURjBn0xxK
RFHY6nHJ48YWx/nSwNOqfD4B8/+aTQChARJ11QbPpQNkegaunOL+da4Wgy9gT3punig66nQML37H
zrmI3uBpKCoIoGCVFMOScJ4woPJRwsH5e5zj0ucoRnRDOKtvBQ8uJ92ojAdym3AjXqcSiu0pY4a9
1M4+DPxQcU29ZKUQrygcrGwNRAOb5nux3fM/kM0FOFfgfWbqYo52oJZ9EB2s/AQI46KE/jYKOwd6
C5WdbzYYerKNyzk837Ki3YdMgvQCiCh3x/URDcMm60JwlwGo4HceVUi3AIOwtp9n3+SqxupZ03g9
szhU/5iHEJ+SSK6vp896+lxVdbufe5j2EB+uXv3vUc6O5dmoR9LvtAwmRGYDS7LljLnMaxI1kAIa
waEEuHC2xOAkDc/NJMQ3+XqwkE3ZoReuZ0F4Qi5Xvp5JWvZiivLW+yVqybAUa31gB/vpr/tRPIZo
+/ZTTtdaxdN7wJPAOXwXFyIeBzrVKEPG4IqFjSqq3XtXcKwFlf411batgjWn6RG05YO/SYJ6bVaC
hLLMqMKwG6X+coJuOJKltYuPNTM3ZqDI60PPEzT+C10TeFvVxc6UXu4kspV/VRQMtnf04W67PWFc
k276F8mSbwxWmWxXrZ85JJvDkpJwcaFTikzhuzSzpbRCioKKpXNYP1oUl8ogrY0ok8J72fZWFPGo
rCMmwJlLJtXcqNOZB+K81g1havU+IXN3BPwLNwy4ZDvpOMsOIMQhRXOPJ9LAJyY9bQQTKN18BG+H
SVDD9VcsZ7QI07vM8JsnMYqsTFe7VHwXUFmqBARovEU4sXLpL/i3jr5H3+0Q5HcjRl3C+GdLYVGN
MPWWYa+K7PuW0KeG9QCvCzvLCbHrx1RjopLJZJGa+Mq5QJCtMR1IHq1+Bdry4FB+qUwQo6xx/Bdz
5qa7j3uxsS7944kqO2fRd4rOnFrAcxc12sg+JiD36qeQZ0svrDghTYENTHD7nDO6V7sgVg9MoXfh
UA7RnXGNQsnLO99FdM4JOp+PXhwZP7j+HfHwjCVzbMOTwtUIKCz8xW1E/SGpo8dPK0nfsh+Ukwq9
UEVF8Lj8kK7EpYB3jj6OhUFLoF0N9u4ksWt582oyAYm9MCWraueiqpFI9gmEIpu5l9D97cpa1NeZ
bf/SiMm6KR+dDIUY8lVsCDv2mNl9cLgkTOOZSWVCG+n4p14sotlOmBq9zQOIJJIPU5kf0BCvDDwR
bhCYZTlCOJZWK8Yj5Kh30sjOnqCpbNLQLVUCGUh7vt4I5Nov5LzFDrtCA7hspnZpk6CdNkwHPTxz
7KyHFWIRtZzkzkYOSar/c9v4BkS/P3VYN5f+i/FBhh+qJZzbLiNj356GsnFMPuFpxFWgzGKosHMT
m7QVRgOAY7PrFSGURCooV7WxopdUNQB+nMaUlrIirrSOLOiql7htuQZbHDHlXRpvDXn4kxmNKfn1
D56K9BAF1PtiGbBv2rZ4mbXgiDfkRFTbT6FKpTibKs+Ev9/Th2+NKYXxijdqvW35m/spoeVY75/s
B4YqZIAc/50w1vLM8dcRtKk+/RX3c/SHAS5ZLdprkKc0WupcCGJImc32VgtMP2/rxVDc0usrhQx2
Wax3O/Ogj7RQh//YLwe4GCBdQv5tbcMGXsXgzowiqHKzuXivI6ftdOd8C87cvDoRRwhty8/axHeX
I/tYpKdufjnrCa9c6gZ4wag7IWDTb/+H59ENTJpuLN5EZyqDzsu64+zqRr5Y6TQujL4xBF6FNEbJ
wdVcaUoMaBJ01Tqy4AM2ANExmOWGO/5IBaWwwiNkxtRcyz3usZn97hO93LKEYVrZYvMg06f+CxLn
yUtOlbo2JRGSnQ9j+AB7yjmo9ffms5VAJw0BpCKzpVwsX/fggkATYriDihew1/2+Y4pMjjhNeaGK
3W9hw1F4ScT5yDbOljAdJSApTnGMg8z3sW7SbXc+/oXq0fS/BgjZtyxjY492z8hvQ9eBar3Hv+dn
5q/SEIjK0BWvcKBe6FN0fgPCd9PmTO92HVOOMBaIAGHxnZ0fOoXMt0wzH+8SJjnK/ryI4qiZtjw6
vRlSIpI0jXi66tGeVM71iDrZ3hQDGQoEr9GGhRwamqv1nhdRxY3nsMubJh2pvNOk1OgSsBa85k1b
ftIpjpGL/ZoXMvn3KqbfgY8Bm7feu3W7pBxa/hadLZECEHddWhv1Z4WmGoXaMrkSeBcwXAsyF26Y
FCxcC3EViT8eokyYKg/mK8q6ByP+kynC0gBWgMQaUb2IbQLIfEneT+Up29Uv8Yv5bB82RW5THzKG
13r7lVU81peanjJTsrAEtZniWYCoST2EhM0AJgPRcIBDA/sgBfvi3+k0ulEcri/wF+c8LPn/8/th
aJLceLqWvd3vDoyn0DdWrHznrv1vk00GGj2MEDvQtpgsTz6NW3vwsb/BO62d+ypXepacTvtxypvw
vqxtp9Lch4Hm2uuDyP2TyexA9WODbEo9XC7AMnt46MZVH+Ro8Azk/vzbdQpOGhtgksvmPqUU/Z/z
U6yeLjQKelRCRrDh+SregsW05aV7zo5QEkbcD7ESj/zU+fRrDd46hWudoK2dT9dVKkpU8mhGgN5n
tFfsrDgvGd3ydyKaxD4QDaVceZ7DhhO5jJow5NJ/6zJ2714+iTTuVR5Q+6AKwrmcjLheyuIntgv2
tZGNUvZE77a1KopSP/OClsuOx8VB59UzCulwbpmmBdW3tao/DlNQnNAJHdSKrt9aCptJIm1FFoXs
cXMHxMLAskI2/wT6idVSrZ2y7AXRCt8tCF+puW5o6zwS1c/PpraMD00BcNpPaEEUDlEZldxs/TqT
WBGjCfqmUwICraDL0kzGcHt86iptsFAkb9XYnmeT8hKGjOMED6Z1VVlwMn543d/6tIpbHvlnpf7l
mwFr0aOfjNVhvxFKTmDuKWRpMNxrU+NxdaYeUEmopJbHu2Ocwvq5r1kJyXN4wKX/Lhroo9DofKj9
0VSdYmr1zPSOVrxnY6PfQ/e+0SF61XpLnXovGwsVrAkGDLgl1opg+8XvjEHZhq6h3V6nsmJkK6b/
xiBMrQx6Ub421x9/vUVXfIxe/S+NKauOCEEri5KVI/Hs1tsLdZAe27yi3uAA9PXM16I9+QdiqlsP
flRizlZdsKe1XS00Yi9TPi4X7RhnnEWSPCxdnT5fIxlyOf9SX7j0eqQ9rGsVWKSh0SuZA2U89dMz
BvvdYPqMhZB7CxqYOK4Djif+nbtXeRMR69CX0VMnNS4mBgeqvHlKLo9arLvwm+AThJ28efzgm2vm
YZtaVVrmfeBcLPHa8SSt2VqXU13iVURqmrNGImlzverwZFTEzO7m3RIsm6UhB07RL4F1RkNYplLK
C/q9Wa6+Yac5oY53rRdbFtpYlJzHM/5cktbMILDReapAS3VvAWC0EyRsBof+0szjn38w+TOG1jH5
aRG0FLxQpMI5yJwBaFirDUWn9LZqILDMy7pIljKxIMSfbUqSUzimb0eRmWkjLAEC9G+9pWbXpuNW
9MqyTwstswlBYRdCQYmBWrkLRjBTTokS00ijBqSyiyyLAuJCy4AfIRtvDAIYYVdyJxdbTTreiL7X
Tkkk94kEZ5zDDiaulEh7v9nMre8Wzxzvur4l/zd2kIucdGhKAmS0ImQpbU3NQYYs+FUmLCwuvfCh
n/EYetzI+DertA5AtFOH6g8nOnPH5BOqh5k63DuXNfVIGY2U5fAp2I403ZL7WvuZh7UsyF0tt6BO
buo7MIXuWDwv2Md8GxH/q3Iuy4nFywWix0+oHgwZiJUlLl7flk7WWpusToINm3rHSa8jg8KLz9ld
FRRc2BeYObAlo56iFlFD8IUJWeborr1c0t08JgIQFeNQJdBmhWCqTt/2/zkx5Z7KfCgQTjCkVufO
ULtwhJA8Z2sKwo3h7rDtGSn/FwQxUrPe1RkfWWaBB5VUW0HX8QmLyc9d3QvZH8FQYc6DM9N+2MAD
HAVw6RYHZx4fQTGgD6MQEZuI99ixtJtXZjEwQJHD5SE9S/skq/E+oWkjYWbsqFSH7wOEexAlYfzy
GCKl5BHMn5iuXD+BnJ6ReeCiM7UU4WUVNgcoJlLRVsYsZUmBHpMXUjeOXPseT6tAJq7MbufchwFz
FHmUNEQ8cA1rXtu2udsujZG+TnfYard8zEOth7SmYfSMgHHD4JPwEN5N7y95q2yDpkdOzIOHXZaE
9FK7tzlDH/ZTBwonrL6U7WMoPD0MB6l+bEABnEHp4fv5+4dKcG19CuRFR8SdDZJ2NGqYY2WivECI
jt+j9bdokzq4GRVRswo/e9bdmXxIT0qZBT9JpI4+us4JR91sRLqmQykrHFRRYfznTHAzcyBrbT0t
jV0q8l/9F6gIB7EFyBIjYd7OnKwzRXJC3tMAgXqxreKSdKFFCketI6zZuPM10vfrO0PDja2pHM7x
1mnNYsbSw04kpewf4+eylrbTvySww/cRnaeAOdh/H/+D0Ok7k/T6aQjFvqGsqfm0NGXmqUaEYIzi
SFbKlWmZrNkVUf6q/S9O/zk5W9LfY6PohitSGUTRG5hk04gwzwsDTowdgycWP/Bd+cg22DBoDH21
Ji/a2+JBfS/HVsajbMELhdhDVwxAjQQ8jjBMp5jVCLUtVo2xnqIurJ0vXB6ICXMJUjYd+a+XiQ6/
yn8xFg90fQL41krFlciuioV5ADh+ElNKLEl3aYX4rWw3osUsR0deXVWJFfVR+UrUdoSMfro0kJxu
6ulFC6/17RnzqBYAYZyqFXRe0zXost17GznARU8zBEi11rH9oudm1eSG7qsxKSrdgzFl8BGf4ITT
COyupcTadw8Lcjdgr+EQqIdEbfX9D8NxabX27J11CE1vrMc8UY7cnbj5WhVLzFKjw5b8rTHaaqE2
VnZPrTAM6SkRvc0EKec96SXFEGNbEmmvHXAi/XQDFjB5CMr6chQ0GzDBuP4PmaQ+Uih65nI7ASG9
PE8HAI/93UqXy16kfJ28QNbzF+Ov3BBN4kxzDZavfAMauxuYM56a+6JFQ/4Jd1Yf6SbxlIgKHjSD
/yYyAAAZRchz6uZLJBWrsls4FJC9BAtPe+vzWCVi5sBAA49TfgfWbK196UKP6T+byTfDfvtXB1MB
sG5cbiU1CsY825r6rVXJtUXZObwRp2Qs3de1Y7JtWYoOvydRSMb12mI12lqYCMRgQ+/X9Oh0GSKo
wcgnpeqo+anuK6mcQXG1Y7LbGWgoFQ0nARn1yOmiLttuaE2iT9aRodCJJSo5+jaiHO9buimRJZKO
KkAE4wPPpBCtyOK0wcdQABhVWEswa4qmHHYbzOHZRH7Wz1PLPersZf7WmYSbaXa+8Ssc0bHeVlbk
RCHtzRBhWf9u9pUNq3dqYWLjC1PiJwfiJxwRR8nXYnT6aEh0c33+9SCI97+9l8nv8yrrmD1qh06O
4GrsmZAF4RzQBQPHrIccU8m2nWvBaQWStTBNULGOlKVVcIdh1Ji0bx5Rldgwh4BBCswuJ7l+uLCD
WF7rtFfqrzJslUHpeKtiITHWm9yPtq9FVjWvEmjzFaagQYkz3rTceF8PFTfw9JJuaxYY9x+9d2gY
DGSdM2FndXIM6H2SMMvgf+DjGMjQeyiRnpAzj1AzxXYaX+hV8gKLiihagI4mZDYFSBLCy23JweAa
SUWXuvQr27PEOCHXem22iI3GRGu3r8fONdAj8FECYIh40iDk63vHd+1E1BKOGRH6Bkqh6o94Ry80
+YIiiv5qnF6FRCLN5ANf2Xq57kbXLl1fAYRWB5YQFI44MiZw7KypojbiU1XBDyekRj4164n9JZZo
70rtoZIv1EEi6PZQmhMpzqM9tlGwpvoXqNAam1Nqast52nNF9PtDs1pxrRzzTXvVMmDW9pUy/vq8
WUrwLTEK7m4gS5m8K453xDLbEyah3YgZxMf+413h02b6aBH71aWiUy5CHjR6WBi7Mh33fnCqlBSQ
I6Dyn5F9QLQM/fxfui73SZeJbyrbuGT0mI7t0YrNd/2cC5CqMpfzkcQz1nuoJcK8mpVIXL5+CMW5
djH0C1dHHH/OP2KiMJUndTqoU9qaMqKaLFF3NmFV64Nw8kCqDcKedAvabGbLGvXbgcPWTdV7iPBg
gR9A640joAXmbUpd63Tg6ZqMVsOr3veNOTmre0HcfaRg+3mVeOcHenRoVqVVJvSldK1Ao6cq5t6y
VWdnQ503qJoo2zmmGEq1RKNjWiN5b+V4DwIED1I++B8jWf2uAkwe9z4MRcgiUptjPPrHtryK/vMd
PQ/4KpY4gRto/REtUUARNynGC2zzixYIBHQukD9mfRGvXTVsvEbHkK1DGfeqSVTMpNFO6ZB4V0XB
99UYjCNuDo//u3phTGtqHCOSyY6wQm6TQ/MHlXOGP5Cf4ogGmpJF/7cSuF4m4HToqjA3IaPn9EIw
g1JQPGKNVfiyGZEfA2MTL5zC9L4/A6CHJ2yl6HK18xDvPc7+T3DghYspD8exftKzE7XRN7zvwIct
xYFitVD9/oXvJM3SaPLg7HrLkv7Z0VmtCfKLNLiKbo77HIAOhhRZEPqs+21O/IEB0/27LQQJh7CV
SDSW0Ge2R+NQ2fUL4h6WGzNEGdS7lD+984VVaoDzTH1xYb2Nh2ifEkSluhsCCp0DeSGThVdnOWD9
bHB7dotf+sitLBaL9PUhueiK51Vb7labdlWmyMVXozZezk+U2noVTxAT5ENl4KlcOvBZ2Zb9TrGt
JEV4uZ7U8OZ4lZwhoh8eR3prWYj+QENHb86LeDy4jmTBGtgNXv1nraK1tGMaiFRMqc5QwFKjD2Su
3WrDECURwJPpRwkD/gLu2snEpU9QfgA/AojBuxwzKD2RhD495LCpNrEGQo93165p/LG6h90fqXV+
eKU9ivgBLi4SzSr7KMQ+dkRtO2FntUlnSSfg/65n0J+TVVKMwwk5Krkg5IMbzJCawgnku0xPx0ss
h1pCZEovcsurMe1lwkseeBfg/aKO5SzH+nBR0PY9te5/tU8rUl5MonDF59yr79OdVfcuRa8KbBGS
kSADQ7MWWdpCGP344VnQr1frYxyjNMS3eSmfJGzBqj2n9xSK5dUmcynY9+i870GpZSjPiCb+Qsp3
+abR3yXaTPMUWKc6cKss8qFEgjANlFKud2Liwv6NA/Aohlyx6REQoyXJy68MRe/kkr8CtgdaomU4
hlHAbDX+d6AM/nVkoEppeKAoFm3+CFih5PtF4M/8INVDpBnk5vIlXM+j7cGXMMG27pfVeTlbBx0c
4K2vuJfFd7j22avSXb2L7+McROxfLiWMRQc79FVgZKh/N0sp8Wzk1QG2gx2RBVUSN3YyqgYSAhoz
1fD0PsFdLse3+uDWP0elcPhA6SZIltb2tloLDJVkdA3EZxc9edwaTwWs+k9tCJ47NqIA6O3nAMJc
UWI9Y/+/TrsGCfx74Jgaif3F7H2vu32dWLj2R6scHm1N50feA4RGAnUIRR2iKyosVg8cjWVP2/Pl
SbCT7dcHQ9NlZBeS4YHuKpdbXOH1EqEf3rRFD1WlCK4S8fgZ9XTjpSUeVfT78kD+WdzgGHU2Ql67
EK0TgJnJK+GjkGY5Zzv2ciSX3UJVDndPsXUUU897J08+v6mqzEX6OnDYvJ5E9l6u5Wfo2/xhRpKZ
XqBF4mBkkuB3bz0rcyza63u5NV/BRlXfafarwG8STRUEr5OZyN6oUaoorUr77wqZJrqDJi/gyR4e
4DztEhLDaDKfpsZkocOrMyEiPyGFJaT2holBew5mNMtg/0mr5uZfJo45Kmu7P6iUf5UaGAbWpHVH
wj9E1jUx+/7IQIYACEHO7A5lF80rYWH7lQLk+znWidrN56hsJWzmPTo83CDIn6GRZ20sD5loSzNS
/dbGNMQ12L1S4y+CHJjQscD3X5tzuQuKwxTwKEDcPwUZQbpZEstSGmejmztDwJdoUgcndau7hyuq
MY7gTMWx5hIluF4xQL74fIq1RI0n32SKf3mhmudY5lioYNJZ6wKqL91dbO66Cs5WjY5rx2AGVw+0
H1UCV8jLodCn+QuGd+t6MPNW44UZlrcM+TOldvVqK6sgp1PzpeSKzqjX4V3rwSpKYfujhlgMnMLb
eshlmSJkYGz7bFREoS27mm3/pvk6sinys+p4u6vWnnasCzAMCVdUYAqcx2TgEJlG7yAQsEd598iU
nqhJHEY279p8EdUh30MmEAKkMAsyrIU3Kt5/1bpIgPrd8ST7a6t6pAI8q5YLZmgyy91itJUMdH+9
dAudOoH501nh91k7vqYzGevQjqDWgiA31dVvo68Si3/cjew4UdDMysmWi+8UyLgbXiJV1zFsSD/o
p2GJqBdSyU1BUH78SRR3QsBFk47/AVIY/JTK2VyR5lCga1Zf3DJ98woDWO4Afw2nGySrI52NkSHs
r7ZK/GbSQQqrB9RXio3BFcRYtn2SNGXRRMz794Om1P08XeP8KWBoo1Z+bC3K/o4giCmykum/D7XK
k6y61WA58EOVm9U2UYCaaHl9nPpZg7kJoL/SXgslS0oVYmYv3cntiucn4fgl4iOhwmI8H+11VKxa
Zoiu2sRpC/ZQLVagg+YZ+Jwp2ab5PJN9RCPbLXL8pluMHvW/fs8zKVsKvmTourJJuRGqoXiZDP0C
gXLwxcPPH1geivSHr4+cKqqriqU9A8Rod2gjZpCkWmmtszphaYOxmuWilI5Y5bZxc/6bfMBr2WO2
67DNTLPUVtTWkxfcJeTIMGwCdsRsYpn2iV9aulyAcjW9k7ubI3UUL1oIOgT1Tj12RAJqpHqKa0Qf
WKo8kc0t8dPbhWgXT4SF821FPLzhdDf9sGO7RznRvtRIW4L8dvAEsyiX0lV6J9YcUlDaBgZlYSHC
6Wp9sk9G6JIu6853LEC954KzadmRBvu0DlUarABU29jOSf7x1p40E8lusRLz4FDUbK78SAiMUwTL
JNSxdAdj3VOoHIyX/Gcl1DOrE7lnkLpJjwKqdoavZXNhFfTlUBzT1JitUPZuucgqbEBoeoNcI9nI
73VQzcEf1C8fEEpGFdvtESOFjefJ8w02lzoGgDgnmuX5GepgAoIcjveorAWWO6hVj6/ItvhLKHCJ
XnKKgUvIq2fBhhOOKdkUKm/ZzrA6mJNy2zOsbamM8+mVNpGtK3VUg2RmAXapBRsxi8+xOrYcuWjo
My5N8zf259ux5l5u1a8/msFCUNLqjBAyaOXRI10EOt8DG/UgAo8xjt5UtbmFKVrEtEVLOPnqfc2D
wC6YJhPUU4ZDsxALodPgK4Any5Mes03we2CLnP9awAe+Vz40VPbR8ioGo4EOk4sRaSw0GuG1fD2+
E+sfG1ZStpkLtJ7VU9sGblTWskqbrZ5JRm1JvyPaeJVj8HrL7VNwtfoDfzHLVadzOm2o4QqA9rQo
Ln6Saf7FStqCv22DV5Tgw5NZLBk6KJ/vWftYyeIVkcq8U5VFqfBAByvrRu5fCpYhYIcaklxlrIsr
r9vEYmbne5PEAW4eFOZdSFFjLtDqIDs/wSOZ98GE9Ua/RLrklMULP+H8kFKcuorItjfYaspI+MiF
zcyfqDG2exHsYi+9Y91Ubqm0A7uypA5ILa5HzKQQ64KC24pYdwVPhcqUFo649fUeRZPwsQtyR9id
61kKAEi2HYlTwXhDBMfLsHixonJvzDb901PikXLJX1NvoZ14QT1LIy7C5W2LtZ6QcypljBmV/ZNL
6FRoNjNVD6/XeX/2/XeCCuSm3y9zWEnWFSjYABBq4YCkA7Y1QLMDNMMFmyCBuuJEf92+zge/Sk96
AsnbgKmHPJhE1QJTcktTFAGOH6k0jIyaykKe7DZ3xcpc8O93W6gQjyOIiRzjAreL+FvZCAMXrFIK
mo81on+e72qpQEgk8Ft5Z/EKLZSC3a0JVEUu9UIskgn7qErHWGdAI5i+BXTVbAF8t1vnPGAimwsF
3Y5zCQTfmhIV1TBW4qaP5BGGzoKhMtQjnxcJFTj8aocpjUyEKcD4n26yQgdwEzVQ+sYBDZt2LzO6
T4rwjf/Tl/99EWBjpvPntZBiaMYIt4ER5sz7ZRUEL355KbjqfCgCVrtGxHPm4DtsNQDtP1FRNSg9
5lq7i/yN1WaxNztkcjCcPkZqOpNuU28WGiq8d0G/FU4xZ26O+Rx8lFISvL6L3BqyeXPLiFFvhgJN
H6TTdXzHJgT+C9mY7YpTAa5kqTBm3htoCoit8wyUsyZY9JUGSXCNff3A3H+Y/DcnLy1YZJKZvtHm
6IMYRy6HR9Pkqy+2rdcnII/mAHFOtHBeAt1hHG92vI+yUcGhsN003QwnTnT/tcWk+Z0HRkJ7pbf9
+OAsWw4tbhgmOKKUa9Jq6MP6CJz63qwJqBGL3rW3VNY9oou8nA4wsTNNWHrWY1cqFRkT4MVgUquH
rXPntyP2HcaL5TjGSmHkbGlhZvc2tMdaxhnMMdvRN008IpkV9hGI2Had2dik4FRMlsW7TsX7FdPA
qEL80Wcb2s7zDRi0FkLJh9JRXas8OIT5RXhFYGaTHM3dqaUm5tcGR3BTxHlli4hplcnbplJbzznS
kQ2ov3tTada7wC2RJGDDs8LWwVw1lKZeV6VrNxNIUv9rDCRUjCOFyEZ39Ioxk9yTHpXPXrqM9VhZ
Xfb5PupX7aps0Wti3iiMy1jxSSAoW7N9zCWg8Q3+R2cWkHvCa7g283TsG+394JBe8LTqbxg2IeTG
U8+ioj06d1zWCJGX0xrBVIL/Vl3pL3LASXEU7ju5dJczPJNL+GYKzI7/sK6XZzRfavTXXlQ69O6l
ZUOcOfiSianHrMs7KdMRebdBWvq8/uBIcFzU7anAe0mvPMMc0iKygWzcfdccaBU52cOfxJpDn2Dh
zlyUWPryMjxKtBRbsVAVpIbYZdi7ClYAtYADl2p2EFhTRAqz7xGKrSCfLTkodaaRWWmhd3wGgigS
/wy5bduDxr9qgzPV5sg7uTByGuPP5Jmpa39sQMZe0l9F+2Rgf94iYAJRrJT6rM+fchEn4Zycpmx4
K4/3Y4lDAWuKXwI5dx/vAvD2CwjSx/nFcVgdV3tmuxe+bUVmraCn9HKppceCdoGRV5moJfvtQ8Hz
Trddn9dhMDsDcUjALpUn1byRx98QH/M+kryyR/Tlgf0/lYX+nPJc6sci45Tnuchppi9A6gzg5Sxg
zGKZYCgesQmKj1IYut4eLxFhIVp+aDXnAb7BBHtbwH2HGnO/eJJPyQrBEcULPp2zvNyzDQveomMl
WncEstn8K3YARSPrDIHf8ZH4gg3gL8KJLBw6+QFjHjbTu7xMdvBQaw+NINYNzIc8cGzjFmlndQe1
jL36SkFD2CEv9OGISRbUg1qN+6FjT8nnzcMjjXZsHt29U9qNT/Uiqc4mXJAl4Tzl1S3jk6fT869U
5q1cZiYbNceXg3WhfhkdO518EYgHvn2hnIEQuMhqrHkko7wAf9hw1mhSipOSIco9uabFZiPvAcbO
/muw1NvgIH2CyuXjLc1ZBhV4Qgl9ff6zbJbFrS1nRTN7vfjpCJFDM8JA77YxNRrWFT7xA5arPkGq
TfKjeswR7ZnjIqrBSq4qwVQQrmbVrXbfSnYUZlwltWhqcYJXYgl8VzOYsjBMrf5FHAdSm4Rkzsc6
+2ny08o5Ch+eF9pz7ij5faDyl3+wBLkXrHi6tRu7RZ7yclrc+WZk2OKt+MHGP61jrHPg0vudYgUt
/MPebnRjesAw1m7EyNMgmLigdAXHF1t/9OlNENYX2JrW8t2f8MMeyHOf+jVGvC5PSBFVjAHzHtCt
LVh07ODy1oxsr2qFmQCv8hx+l6VGxGWpGnytoNsSU+4oWgs8UpomBQzy2ioaLbNXSxd4gUw8w44R
WtMbAKvWELpwdvJT/ekAOJPwAIRRh89nbCB900ova94AzVnWpuE5sH3mT8KBEj6Zmgk1kPTaDEDa
IG0UN21OVjNSomx3XRrvmbTIM6Tx1btwiczNIDLZYN2IXqCIjr5iDtdxTZ0K0IPf8Ef7Zm71aMTS
TE72/hcN4XgjrOyXv1uu6gyDIC0JLCDpY7MUjmCLOtkBNWM87qHv1ykuPxeJc6ZRGF32YzJgK1Wy
2Vq0r90zkpKFHtPtRotzXdVmC1zZc+GtVmM70aeO1IJWzYv2S5EwCciTOs2UgWTHvm2hQfVQJAk/
+mPw+KkYAQIyqE9JRwuDEggrwbS2HiNP9w8XiaxewuccJcgYZz1v0D7B8uZXRrtFFiEZtbFti9W9
vRTR9UTeWVxcu9eHbLXVkOqtiBd1xhnf635eNPy1iulH99PRbh2SDuOsJz25k14Qv4mhQaNQahby
ICeoVJoYMvfI21eHwKIIseYlT8Lyhy3eenYq5G53SuQ2e1/wintFwre7mptn2V0hj/HJIBmfJ9qt
+bE3NnHVpY0hFi9c2LKboOKNP9+GBvnwVRYn3KA86YsidBbtpyJ1qmIkbJYjIGLMFk/mDOs6kLiA
Rg==
`protect end_protected
