`timescale 1 ps / 1 ps

module altera_highspeed_rs_enc_lagr_poly(
     lagrange_poly
);

    output [32-1:0][32-1:0][8-1:0] lagrange_poly;

    wire [32-1:0][32-1:0][8-1:0] T;

    assign T[0][0] = 254; assign T[0][1] = 60; assign T[0][2] = 161; assign T[0][3] = 131; assign T[0][4] = 186; assign T[0][5] = 216; assign T[0][6] = 247; assign T[0][7] = 217; assign T[0][8] = 102; assign T[0][9] = 75; assign T[0][10] = 248; assign T[0][11] = 124; assign T[0][12] = 116; assign T[0][13] = 22; assign T[0][14] = 139; assign T[0][15] = 1; assign T[0][16] = 22; assign T[0][17] = 87; assign T[0][18] = 115; assign T[0][19] = 146; assign T[0][20] = 72; assign T[0][21] = 100; assign T[0][22] = 72; assign T[0][23] = 21; assign T[0][24] = 240; assign T[0][25] = 196; assign T[0][26] = 215; assign T[0][27] = 14; assign T[0][28] = 68; assign T[0][29] = 21; assign T[0][30] = 197; assign T[0][31] = 68; 
    assign T[1][0] = 68; assign T[1][1] = 197; assign T[1][2] = 115; assign T[1][3] = 203; assign T[1][4] = 23; assign T[1][5] = 77; assign T[1][6] = 19; assign T[1][7] = 47; assign T[1][8] = 122; assign T[1][9] = 160; assign T[1][10] = 103; assign T[1][11] = 132; assign T[1][12] = 218; assign T[1][13] = 165; assign T[1][14] = 67; assign T[1][15] = 100; assign T[1][16] = 102; assign T[1][17] = 148; assign T[1][18] = 92; assign T[1][19] = 166; assign T[1][20] = 1; assign T[1][21] = 0; assign T[1][22] = 142; assign T[1][23] = 25; assign T[1][24] = 70; assign T[1][25] = 24; assign T[1][26] = 20; assign T[1][27] = 109; assign T[1][28] = 178; assign T[1][29] = 211; assign T[1][30] = 11; assign T[1][31] = 237; 
    assign T[2][0] = 31; assign T[2][1] = 149; assign T[2][2] = 216; assign T[2][3] = 80; assign T[2][4] = 95; assign T[2][5] = 120; assign T[2][6] = 111; assign T[2][7] = 160; assign T[2][8] = 244; assign T[2][9] = 74; assign T[2][10] = 84; assign T[2][11] = 132; assign T[2][12] = 57; assign T[2][13] = 239; assign T[2][14] = 72; assign T[2][15] = 145; assign T[2][16] = 90; assign T[2][17] = 91; assign T[2][18] = 179; assign T[2][19] = 219; assign T[2][20] = 140; assign T[2][21] = 87; assign T[2][22] = 168; assign T[2][23] = 205; assign T[2][24] = 70; assign T[2][25] = 195; assign T[2][26] = 204; assign T[2][27] = 69; assign T[2][28] = 136; assign T[2][29] = 209; assign T[2][30] = 30; assign T[2][31] = 23; 
    assign T[3][0] = 194; assign T[3][1] = 192; assign T[3][2] = 240; assign T[3][3] = 227; assign T[3][4] = 155; assign T[3][5] = 40; assign T[3][6] = 67; assign T[3][7] = 95; assign T[3][8] = 122; assign T[3][9] = 229; assign T[3][10] = 106; assign T[3][11] = 217; assign T[3][12] = 61; assign T[3][13] = 245; assign T[3][14] = 213; assign T[3][15] = 1; assign T[3][16] = 125; assign T[3][17] = 251; assign T[3][18] = 40; assign T[3][19] = 156; assign T[3][20] = 130; assign T[3][21] = 1; assign T[3][22] = 251; assign T[3][23] = 105; assign T[3][24] = 242; assign T[3][25] = 143; assign T[3][26] = 110; assign T[3][27] = 203; assign T[3][28] = 191; assign T[3][29] = 175; assign T[3][30] = 14; assign T[3][31] = 107; 
    assign T[4][0] = 213; assign T[4][1] = 221; assign T[4][2] = 62; assign T[4][3] = 176; assign T[4][4] = 2; assign T[4][5] = 117; assign T[4][6] = 185; assign T[4][7] = 83; assign T[4][8] = 133; assign T[4][9] = 232; assign T[4][10] = 172; assign T[4][11] = 97; assign T[4][12] = 187; assign T[4][13] = 40; assign T[4][14] = 174; assign T[4][15] = 75; assign T[4][16] = 248; assign T[4][17] = 161; assign T[4][18] = 231; assign T[4][19] = 139; assign T[4][20] = 19; assign T[4][21] = 36; assign T[4][22] = 21; assign T[4][23] = 173; assign T[4][24] = 16; assign T[4][25] = 254; assign T[4][26] = 208; assign T[4][27] = 156; assign T[4][28] = 244; assign T[4][29] = 162; assign T[4][30] = 124; assign T[4][31] = 255; 
    assign T[5][0] = 118; assign T[5][1] = 233; assign T[5][2] = 146; assign T[5][3] = 136; assign T[5][4] = 159; assign T[5][5] = 59; assign T[5][6] = 56; assign T[5][7] = 171; assign T[5][8] = 146; assign T[5][9] = 88; assign T[5][10] = 22; assign T[5][11] = 13; assign T[5][12] = 163; assign T[5][13] = 94; assign T[5][14] = 0; assign T[5][15] = 1; assign T[5][16] = 211; assign T[5][17] = 46; assign T[5][18] = 59; assign T[5][19] = 144; assign T[5][20] = 244; assign T[5][21] = 9; assign T[5][22] = 6; assign T[5][23] = 148; assign T[5][24] = 87; assign T[5][25] = 215; assign T[5][26] = 178; assign T[5][27] = 68; assign T[5][28] = 241; assign T[5][29] = 189; assign T[5][30] = 24; assign T[5][31] = 132; 
    assign T[6][0] = 204; assign T[6][1] = 66; assign T[6][2] = 209; assign T[6][3] = 246; assign T[6][4] = 103; assign T[6][5] = 72; assign T[6][6] = 124; assign T[6][7] = 88; assign T[6][8] = 211; assign T[6][9] = 164; assign T[6][10] = 13; assign T[6][11] = 8; assign T[6][12] = 24; assign T[6][13] = 175; assign T[6][14] = 31; assign T[6][15] = 40; assign T[6][16] = 223; assign T[6][17] = 159; assign T[6][18] = 80; assign T[6][19] = 195; assign T[6][20] = 175; assign T[6][21] = 44; assign T[6][22] = 116; assign T[6][23] = 242; assign T[6][24] = 247; assign T[6][25] = 5; assign T[6][26] = 198; assign T[6][27] = 30; assign T[6][28] = 64; assign T[6][29] = 130; assign T[6][30] = 71; assign T[6][31] = 41; 
    assign T[7][0] = 76; assign T[7][1] = 86; assign T[7][2] = 150; assign T[7][3] = 198; assign T[7][4] = 6; assign T[7][5] = 61; assign T[7][6] = 232; assign T[7][7] = 121; assign T[7][8] = 120; assign T[7][9] = 132; assign T[7][10] = 235; assign T[7][11] = 164; assign T[7][12] = 68; assign T[7][13] = 133; assign T[7][14] = 153; assign T[7][15] = 58; assign T[7][16] = 190; assign T[7][17] = 250; assign T[7][18] = 25; assign T[7][19] = 246; assign T[7][20] = 225; assign T[7][21] = 47; assign T[7][22] = 34; assign T[7][23] = 103; assign T[7][24] = 39; assign T[7][25] = 72; assign T[7][26] = 219; assign T[7][27] = 88; assign T[7][28] = 87; assign T[7][29] = 45; assign T[7][30] = 205; assign T[7][31] = 74; 
    assign T[8][0] = 188; assign T[8][1] = 164; assign T[8][2] = 51; assign T[8][3] = 134; assign T[8][4] = 61; assign T[8][5] = 61; assign T[8][6] = 184; assign T[8][7] = 136; assign T[8][8] = 175; assign T[8][9] = 227; assign T[8][10] = 197; assign T[8][11] = 185; assign T[8][12] = 76; assign T[8][13] = 140; assign T[8][14] = 242; assign T[8][15] = 0; assign T[8][16] = 129; assign T[8][17] = 252; assign T[8][18] = 183; assign T[8][19] = 48; assign T[8][20] = 152; assign T[8][21] = 51; assign T[8][22] = 228; assign T[8][23] = 103; assign T[8][24] = 13; assign T[8][25] = 56; assign T[8][26] = 180; assign T[8][27] = 61; assign T[8][28] = 24; assign T[8][29] = 245; assign T[8][30] = 170; assign T[8][31] = 182; 
    assign T[9][0] = 164; assign T[9][1] = 1; assign T[9][2] = 121; assign T[9][3] = 95; assign T[9][4] = 79; assign T[9][5] = 177; assign T[9][6] = 18; assign T[9][7] = 174; assign T[9][8] = 56; assign T[9][9] = 114; assign T[9][10] = 109; assign T[9][11] = 175; assign T[9][12] = 161; assign T[9][13] = 45; assign T[9][14] = 140; assign T[9][15] = 114; assign T[9][16] = 52; assign T[9][17] = 2; assign T[9][18] = 67; assign T[9][19] = 180; assign T[9][20] = 140; assign T[9][21] = 245; assign T[9][22] = 21; assign T[9][23] = 85; assign T[9][24] = 225; assign T[9][25] = 131; assign T[9][26] = 4; assign T[9][27] = 206; assign T[9][28] = 7; assign T[9][29] = 68; assign T[9][30] = 83; assign T[9][31] = 123; 
    assign T[10][0] = 206; assign T[10][1] = 253; assign T[10][2] = 254; assign T[10][3] = 239; assign T[10][4] = 124; assign T[10][5] = 189; assign T[10][6] = 221; assign T[10][7] = 160; assign T[10][8] = 246; assign T[10][9] = 183; assign T[10][10] = 96; assign T[10][11] = 215; assign T[10][12] = 224; assign T[10][13] = 190; assign T[10][14] = 0; assign T[10][15] = 233; assign T[10][16] = 162; assign T[10][17] = 247; assign T[10][18] = 145; assign T[10][19] = 243; assign T[10][20] = 220; assign T[10][21] = 198; assign T[10][22] = 36; assign T[10][23] = 31; assign T[10][24] = 10; assign T[10][25] = 195; assign T[10][26] = 25; assign T[10][27] = 87; assign T[10][28] = 242; assign T[10][29] = 21; assign T[10][30] = 0; assign T[10][31] = 169; 
    assign T[11][0] = 169; assign T[11][1] = 169; assign T[11][2] = 103; assign T[11][3] = 212; assign T[11][4] = 88; assign T[11][5] = 142; assign T[11][6] = 133; assign T[11][7] = 54; assign T[11][8] = 169; assign T[11][9] = 41; assign T[11][10] = 100; assign T[11][11] = 73; assign T[11][12] = 16; assign T[11][13] = 97; assign T[11][14] = 80; assign T[11][15] = 100; assign T[11][16] = 118; assign T[11][17] = 108; assign T[11][18] = 142; assign T[11][19] = 50; assign T[11][20] = 245; assign T[11][21] = 49; assign T[11][22] = 74; assign T[11][23] = 142; assign T[11][24] = 190; assign T[11][25] = 194; assign T[11][26] = 50; assign T[11][27] = 144; assign T[11][28] = 168; assign T[11][29] = 108; assign T[11][30] = 100; assign T[11][31] = 230; 
    assign T[12][0] = 160; assign T[12][1] = 57; assign T[12][2] = 164; assign T[12][3] = 7; assign T[12][4] = 24; assign T[12][5] = 232; assign T[12][6] = 171; assign T[12][7] = 144; assign T[12][8] = 248; assign T[12][9] = 33; assign T[12][10] = 71; assign T[12][11] = 48; assign T[12][12] = 188; assign T[12][13] = 118; assign T[12][14] = 51; assign T[12][15] = 72; assign T[12][16] = 32; assign T[12][17] = 172; assign T[12][18] = 211; assign T[12][19] = 3; assign T[12][20] = 165; assign T[12][21] = 69; assign T[12][22] = 4; assign T[12][23] = 32; assign T[12][24] = 84; assign T[12][25] = 150; assign T[12][26] = 55; assign T[12][27] = 87; assign T[12][28] = 203; assign T[12][29] = 237; assign T[12][30] = 21; assign T[12][31] = 231; 
    assign T[13][0] = 80; assign T[13][1] = 243; assign T[13][2] = 235; assign T[13][3] = 72; assign T[13][4] = 201; assign T[13][5] = 38; assign T[13][6] = 152; assign T[13][7] = 201; assign T[13][8] = 241; assign T[13][9] = 199; assign T[13][10] = 132; assign T[13][11] = 248; assign T[13][12] = 154; assign T[13][13] = 63; assign T[13][14] = 213; assign T[13][15] = 13; assign T[13][16] = 65; assign T[13][17] = 126; assign T[13][18] = 120; assign T[13][19] = 30; assign T[13][20] = 176; assign T[13][21] = 41; assign T[13][22] = 137; assign T[13][23] = 133; assign T[13][24] = 213; assign T[13][25] = 205; assign T[13][26] = 101; assign T[13][27] = 12; assign T[13][28] = 27; assign T[13][29] = 26; assign T[13][30] = 210; assign T[13][31] = 231; 
    assign T[14][0] = 60; assign T[14][1] = 252; assign T[14][2] = 76; assign T[14][3] = 219; assign T[14][4] = 55; assign T[14][5] = 0; assign T[14][6] = 105; assign T[14][7] = 125; assign T[14][8] = 208; assign T[14][9] = 241; assign T[14][10] = 0; assign T[14][11] = 23; assign T[14][12] = 255; assign T[14][13] = 98; assign T[14][14] = 137; assign T[14][15] = 11; assign T[14][16] = 213; assign T[14][17] = 194; assign T[14][18] = 209; assign T[14][19] = 81; assign T[14][20] = 247; assign T[14][21] = 81; assign T[14][22] = 72; assign T[14][23] = 184; assign T[14][24] = 112; assign T[14][25] = 71; assign T[14][26] = 30; assign T[14][27] = 8; assign T[14][28] = 252; assign T[14][29] = 180; assign T[14][30] = 239; assign T[14][31] = 26; 
    assign T[15][0] = 59; assign T[15][1] = 156; assign T[15][2] = 235; assign T[15][3] = 193; assign T[15][4] = 14; assign T[15][5] = 108; assign T[15][6] = 201; assign T[15][7] = 162; assign T[15][8] = 0; assign T[15][9] = 5; assign T[15][10] = 124; assign T[15][11] = 106; assign T[15][12] = 159; assign T[15][13] = 57; assign T[15][14] = 29; assign T[15][15] = 149; assign T[15][16] = 52; assign T[15][17] = 170; assign T[15][18] = 75; assign T[15][19] = 176; assign T[15][20] = 175; assign T[15][21] = 75; assign T[15][22] = 94; assign T[15][23] = 94; assign T[15][24] = 152; assign T[15][25] = 37; assign T[15][26] = 234; assign T[15][27] = 5; assign T[15][28] = 179; assign T[15][29] = 200; assign T[15][30] = 181; assign T[15][31] = 164; 
    assign T[16][0] = 23; assign T[16][1] = 207; assign T[16][2] = 62; assign T[16][3] = 105; assign T[16][4] = 209; assign T[16][5] = 68; assign T[16][6] = 214; assign T[16][7] = 156; assign T[16][8] = 186; assign T[16][9] = 6; assign T[16][10] = 13; assign T[16][11] = 207; assign T[16][12] = 26; assign T[16][13] = 232; assign T[16][14] = 166; assign T[16][15] = 92; assign T[16][16] = 171; assign T[16][17] = 72; assign T[16][18] = 177; assign T[16][19] = 112; assign T[16][20] = 145; assign T[16][21] = 162; assign T[16][22] = 31; assign T[16][23] = 0; assign T[16][24] = 89; assign T[16][25] = 27; assign T[16][26] = 87; assign T[16][27] = 104; assign T[16][28] = 219; assign T[16][29] = 231; assign T[16][30] = 26; assign T[16][31] = 115; 
    assign T[17][0] = 13; assign T[17][1] = 196; assign T[17][2] = 121; assign T[17][3] = 137; assign T[17][4] = 109; assign T[17][5] = 255; assign T[17][6] = 97; assign T[17][7] = 22; assign T[17][8] = 33; assign T[17][9] = 56; assign T[17][10] = 73; assign T[17][11] = 77; assign T[17][12] = 223; assign T[17][13] = 205; assign T[17][14] = 42; assign T[17][15] = 56; assign T[17][16] = 216; assign T[17][17] = 93; assign T[17][18] = 109; assign T[17][19] = 226; assign T[17][20] = 45; assign T[17][21] = 0; assign T[17][22] = 2; assign T[17][23] = 115; assign T[17][24] = 29; assign T[17][25] = 35; assign T[17][26] = 0; assign T[17][27] = 129; assign T[17][28] = 202; assign T[17][29] = 79; assign T[17][30] = 4; assign T[17][31] = 169; 
    assign T[18][0] = 134; assign T[18][1] = 159; assign T[18][2] = 111; assign T[18][3] = 246; assign T[18][4] = 227; assign T[18][5] = 174; assign T[18][6] = 134; assign T[18][7] = 242; assign T[18][8] = 146; assign T[18][9] = 153; assign T[18][10] = 103; assign T[18][11] = 241; assign T[18][12] = 247; assign T[18][13] = 224; assign T[18][14] = 64; assign T[18][15] = 142; assign T[18][16] = 79; assign T[18][17] = 183; assign T[18][18] = 79; assign T[18][19] = 214; assign T[18][20] = 143; assign T[18][21] = 152; assign T[18][22] = 86; assign T[18][23] = 250; assign T[18][24] = 222; assign T[18][25] = 3; assign T[18][26] = 131; assign T[18][27] = 18; assign T[18][28] = 21; assign T[18][29] = 147; assign T[18][30] = 177; assign T[18][31] = 92; 
    assign T[19][0] = 199; assign T[19][1] = 41; assign T[19][2] = 91; assign T[19][3] = 150; assign T[19][4] = 68; assign T[19][5] = 194; assign T[19][6] = 192; assign T[19][7] = 43; assign T[19][8] = 140; assign T[19][9] = 38; assign T[19][10] = 224; assign T[19][11] = 66; assign T[19][12] = 28; assign T[19][13] = 72; assign T[19][14] = 120; assign T[19][15] = 127; assign T[19][16] = 234; assign T[19][17] = 77; assign T[19][18] = 103; assign T[19][19] = 48; assign T[19][20] = 178; assign T[19][21] = 164; assign T[19][22] = 8; assign T[19][23] = 167; assign T[19][24] = 96; assign T[19][25] = 167; assign T[19][26] = 128; assign T[19][27] = 27; assign T[19][28] = 184; assign T[19][29] = 20; assign T[19][30] = 6; assign T[19][31] = 170; 
    assign T[20][0] = 195; assign T[20][1] = 172; assign T[20][2] = 250; assign T[20][3] = 104; assign T[20][4] = 115; assign T[20][5] = 226; assign T[20][6] = 130; assign T[20][7] = 115; assign T[20][8] = 222; assign T[20][9] = 47; assign T[20][10] = 98; assign T[20][11] = 56; assign T[20][12] = 109; assign T[20][13] = 191; assign T[20][14] = 204; assign T[20][15] = 138; assign T[20][16] = 116; assign T[20][17] = 182; assign T[20][18] = 137; assign T[20][19] = 203; assign T[20][20] = 67; assign T[20][21] = 103; assign T[20][22] = 192; assign T[20][23] = 125; assign T[20][24] = 188; assign T[20][25] = 241; assign T[20][26] = 19; assign T[20][27] = 36; assign T[20][28] = 54; assign T[20][29] = 157; assign T[20][30] = 6; assign T[20][31] = 108; 
    assign T[21][0] = 89; assign T[21][1] = 0; assign T[21][2] = 57; assign T[21][3] = 100; assign T[21][4] = 132; assign T[21][5] = 31; assign T[21][6] = 26; assign T[21][7] = 198; assign T[21][8] = 100; assign T[21][9] = 117; assign T[21][10] = 149; assign T[21][11] = 227; assign T[21][12] = 65; assign T[21][13] = 91; assign T[21][14] = 133; assign T[21][15] = 137; assign T[21][16] = 240; assign T[21][17] = 0; assign T[21][18] = 91; assign T[21][19] = 14; assign T[21][20] = 169; assign T[21][21] = 86; assign T[21][22] = 111; assign T[21][23] = 193; assign T[21][24] = 170; assign T[21][25] = 19; assign T[21][26] = 84; assign T[21][27] = 199; assign T[21][28] = 220; assign T[21][29] = 48; assign T[21][30] = 233; assign T[21][31] = 233; 
    assign T[22][0] = 232; assign T[22][1] = 19; assign T[22][2] = 218; assign T[22][3] = 14; assign T[22][4] = 231; assign T[22][5] = 200; assign T[22][6] = 114; assign T[22][7] = 69; assign T[22][8] = 216; assign T[22][9] = 178; assign T[22][10] = 38; assign T[22][11] = 186; assign T[22][12] = 173; assign T[22][13] = 238; assign T[22][14] = 179; assign T[22][15] = 233; assign T[22][16] = 29; assign T[22][17] = 102; assign T[22][18] = 95; assign T[22][19] = 120; assign T[22][20] = 231; assign T[22][21] = 177; assign T[22][22] = 60; assign T[22][23] = 91; assign T[22][24] = 5; assign T[22][25] = 40; assign T[22][26] = 66; assign T[22][27] = 183; assign T[22][28] = 160; assign T[22][29] = 123; assign T[22][30] = 149; assign T[22][31] = 35; 
    assign T[23][0] = 83; assign T[23][1] = 243; assign T[23][2] = 12; assign T[23][3] = 70; assign T[23][4] = 155; assign T[23][5] = 243; assign T[23][6] = 133; assign T[23][7] = 1; assign T[23][8] = 244; assign T[23][9] = 233; assign T[23][10] = 196; assign T[23][11] = 238; assign T[23][12] = 3; assign T[23][13] = 197; assign T[23][14] = 68; assign T[23][15] = 38; assign T[23][16] = 0; assign T[23][17] = 80; assign T[23][18] = 62; assign T[23][19] = 5; assign T[23][20] = 161; assign T[23][21] = 226; assign T[23][22] = 237; assign T[23][23] = 128; assign T[23][24] = 139; assign T[23][25] = 235; assign T[23][26] = 193; assign T[23][27] = 19; assign T[23][28] = 189; assign T[23][29] = 13; assign T[23][30] = 175; assign T[23][31] = 125; 
    assign T[24][0] = 229; assign T[24][1] = 31; assign T[24][2] = 254; assign T[24][3] = 61; assign T[24][4] = 54; assign T[24][5] = 57; assign T[24][6] = 123; assign T[24][7] = 224; assign T[24][8] = 54; assign T[24][9] = 162; assign T[24][10] = 154; assign T[24][11] = 169; assign T[24][12] = 165; assign T[24][13] = 219; assign T[24][14] = 141; assign T[24][15] = 176; assign T[24][16] = 114; assign T[24][17] = 196; assign T[24][18] = 121; assign T[24][19] = 114; assign T[24][20] = 179; assign T[24][21] = 72; assign T[24][22] = 17; assign T[24][23] = 128; assign T[24][24] = 103; assign T[24][25] = 109; assign T[24][26] = 95; assign T[24][27] = 177; assign T[24][28] = 25; assign T[24][29] = 171; assign T[24][30] = 110; assign T[24][31] = 166; 
    assign T[25][0] = 119; assign T[25][1] = 199; assign T[25][2] = 6; assign T[25][3] = 95; assign T[25][4] = 136; assign T[25][5] = 230; assign T[25][6] = 38; assign T[25][7] = 63; assign T[25][8] = 248; assign T[25][9] = 158; assign T[25][10] = 231; assign T[25][11] = 191; assign T[25][12] = 108; assign T[25][13] = 186; assign T[25][14] = 45; assign T[25][15] = 192; assign T[25][16] = 43; assign T[25][17] = 131; assign T[25][18] = 28; assign T[25][19] = 17; assign T[25][20] = 238; assign T[25][21] = 62; assign T[25][22] = 133; assign T[25][23] = 96; assign T[25][24] = 183; assign T[25][25] = 2; assign T[25][26] = 231; assign T[25][27] = 87; assign T[25][28] = 69; assign T[25][29] = 171; assign T[25][30] = 51; assign T[25][31] = 211; 
    assign T[26][0] = 160; assign T[26][1] = 126; assign T[26][2] = 155; assign T[26][3] = 216; assign T[26][4] = 82; assign T[26][5] = 72; assign T[26][6] = 57; assign T[26][7] = 42; assign T[26][8] = 239; assign T[26][9] = 123; assign T[26][10] = 187; assign T[26][11] = 210; assign T[26][12] = 3; assign T[26][13] = 42; assign T[26][14] = 118; assign T[26][15] = 181; assign T[26][16] = 149; assign T[26][17] = 0; assign T[26][18] = 130; assign T[26][19] = 98; assign T[26][20] = 198; assign T[26][21] = 135; assign T[26][22] = 22; assign T[26][23] = 59; assign T[26][24] = 62; assign T[26][25] = 52; assign T[26][26] = 54; assign T[26][27] = 168; assign T[26][28] = 215; assign T[26][29] = 87; assign T[26][30] = 108; assign T[26][31] = 226; 
    assign T[27][0] = 189; assign T[27][1] = 45; assign T[27][2] = 231; assign T[27][3] = 188; assign T[27][4] = 17; assign T[27][5] = 42; assign T[27][6] = 163; assign T[27][7] = 245; assign T[27][8] = 25; assign T[27][9] = 10; assign T[27][10] = 13; assign T[27][11] = 237; assign T[27][12] = 80; assign T[27][13] = 236; assign T[27][14] = 202; assign T[27][15] = 226; assign T[27][16] = 204; assign T[27][17] = 104; assign T[27][18] = 50; assign T[27][19] = 25; assign T[27][20] = 77; assign T[27][21] = 135; assign T[27][22] = 24; assign T[27][23] = 62; assign T[27][24] = 209; assign T[27][25] = 22; assign T[27][26] = 229; assign T[27][27] = 199; assign T[27][28] = 202; assign T[27][29] = 229; assign T[27][30] = 61; assign T[27][31] = 85; 
    assign T[28][0] = 74; assign T[28][1] = 118; assign T[28][2] = 125; assign T[28][3] = 234; assign T[28][4] = 190; assign T[28][5] = 22; assign T[28][6] = 159; assign T[28][7] = 221; assign T[28][8] = 45; assign T[28][9] = 99; assign T[28][10] = 146; assign T[28][11] = 210; assign T[28][12] = 102; assign T[28][13] = 31; assign T[28][14] = 29; assign T[28][15] = 88; assign T[28][16] = 138; assign T[28][17] = 182; assign T[28][18] = 79; assign T[28][19] = 68; assign T[28][20] = 50; assign T[28][21] = 104; assign T[28][22] = 167; assign T[28][23] = 251; assign T[28][24] = 148; assign T[28][25] = 212; assign T[28][26] = 172; assign T[28][27] = 67; assign T[28][28] = 6; assign T[28][29] = 146; assign T[28][30] = 137; assign T[28][31] = 240; 
    assign T[29][0] = 34; assign T[29][1] = 152; assign T[29][2] = 188; assign T[29][3] = 139; assign T[29][4] = 47; assign T[29][5] = 14; assign T[29][6] = 4; assign T[29][7] = 105; assign T[29][8] = 207; assign T[29][9] = 91; assign T[29][10] = 52; assign T[29][11] = 174; assign T[29][12] = 157; assign T[29][13] = 108; assign T[29][14] = 132; assign T[29][15] = 37; assign T[29][16] = 170; assign T[29][17] = 49; assign T[29][18] = 66; assign T[29][19] = 35; assign T[29][20] = 4; assign T[29][21] = 122; assign T[29][22] = 91; assign T[29][23] = 142; assign T[29][24] = 70; assign T[29][25] = 201; assign T[29][26] = 58; assign T[29][27] = 86; assign T[29][28] = 171; assign T[29][29] = 225; assign T[29][30] = 207; assign T[29][31] = 168; 
    assign T[30][0] = 208; assign T[30][1] = 7; assign T[30][2] = 232; assign T[30][3] = 189; assign T[30][4] = 1; assign T[30][5] = 84; assign T[30][6] = 254; assign T[30][7] = 60; assign T[30][8] = 65; assign T[30][9] = 69; assign T[30][10] = 0; assign T[30][11] = 230; assign T[30][12] = 231; assign T[30][13] = 122; assign T[30][14] = 26; assign T[30][15] = 191; assign T[30][16] = 28; assign T[30][17] = 101; assign T[30][18] = 92; assign T[30][19] = 159; assign T[30][20] = 117; assign T[30][21] = 239; assign T[30][22] = 23; assign T[30][23] = 152; assign T[30][24] = 231; assign T[30][25] = 108; assign T[30][26] = 226; assign T[30][27] = 70; assign T[30][28] = 151; assign T[30][29] = 76; assign T[30][30] = 221; assign T[30][31] = 73; 
    assign T[31][0] = 129; assign T[31][1] = 68; assign T[31][2] = 225; assign T[31][3] = 90; assign T[31][4] = 214; assign T[31][5] = 3; assign T[31][6] = 128; assign T[31][7] = 204; assign T[31][8] = 183; assign T[31][9] = 121; assign T[31][10] = 85; assign T[31][11] = 85; assign T[31][12] = 159; assign T[31][13] = 117; assign T[31][14] = 180; assign T[31][15] = 53; assign T[31][16] = 143; assign T[31][17] = 244; assign T[31][18] = 56; assign T[31][19] = 200; assign T[31][20] = 38; assign T[31][21] = 44; assign T[31][22] = 152; assign T[31][23] = 165; assign T[31][24] = 204; assign T[31][25] = 247; assign T[31][26] = 172; assign T[31][27] = 108; assign T[31][28] = 57; assign T[31][29] = 50; assign T[31][30] = 219; assign T[31][31] = 213; 
    assign lagrange_poly = T;

endmodule


`timescale 1 ps / 1 ps

module altera_highspeed_rs_enc_alphas(
     alphas
);

    output [255:0][8-1:0] alphas;

    wire [255:0][8-1:0] T;

    assign T[0] = 1; assign T[1] = 2; assign T[2] = 4; assign T[3] = 8; assign T[4] = 16; assign T[5] = 32; assign T[6] = 64; assign T[7] = 128; assign T[8] = 29; assign T[9] = 58; assign T[10] = 116; assign T[11] = 232; assign T[12] = 205; assign T[13] = 135; assign T[14] = 19; assign T[15] = 38; assign T[16] = 76; assign T[17] = 152; assign T[18] = 45; assign T[19] = 90; assign T[20] = 180; assign T[21] = 117; assign T[22] = 234; assign T[23] = 201; assign T[24] = 143; 
    assign T[25] = 3; assign T[26] = 6; assign T[27] = 12; assign T[28] = 24; assign T[29] = 48; assign T[30] = 96; assign T[31] = 192; assign T[32] = 157; assign T[33] = 39; assign T[34] = 78; assign T[35] = 156; assign T[36] = 37; assign T[37] = 74; assign T[38] = 148; assign T[39] = 53; assign T[40] = 106; assign T[41] = 212; assign T[42] = 181; assign T[43] = 119; assign T[44] = 238; assign T[45] = 193; assign T[46] = 159; assign T[47] = 35; assign T[48] = 70; assign T[49] = 140; 
    assign T[50] = 5; assign T[51] = 10; assign T[52] = 20; assign T[53] = 40; assign T[54] = 80; assign T[55] = 160; assign T[56] = 93; assign T[57] = 186; assign T[58] = 105; assign T[59] = 210; assign T[60] = 185; assign T[61] = 111; assign T[62] = 222; assign T[63] = 161; assign T[64] = 95; assign T[65] = 190; assign T[66] = 97; assign T[67] = 194; assign T[68] = 153; assign T[69] = 47; assign T[70] = 94; assign T[71] = 188; assign T[72] = 101; assign T[73] = 202; assign T[74] = 137; 
    assign T[75] = 15; assign T[76] = 30; assign T[77] = 60; assign T[78] = 120; assign T[79] = 240; assign T[80] = 253; assign T[81] = 231; assign T[82] = 211; assign T[83] = 187; assign T[84] = 107; assign T[85] = 214; assign T[86] = 177; assign T[87] = 127; assign T[88] = 254; assign T[89] = 225; assign T[90] = 223; assign T[91] = 163; assign T[92] = 91; assign T[93] = 182; assign T[94] = 113; assign T[95] = 226; assign T[96] = 217; assign T[97] = 175; assign T[98] = 67; assign T[99] = 134; 
    assign T[100] = 17; assign T[101] = 34; assign T[102] = 68; assign T[103] = 136; assign T[104] = 13; assign T[105] = 26; assign T[106] = 52; assign T[107] = 104; assign T[108] = 208; assign T[109] = 189; assign T[110] = 103; assign T[111] = 206; assign T[112] = 129; assign T[113] = 31; assign T[114] = 62; assign T[115] = 124; assign T[116] = 248; assign T[117] = 237; assign T[118] = 199; assign T[119] = 147; assign T[120] = 59; assign T[121] = 118; assign T[122] = 236; assign T[123] = 197; assign T[124] = 151; 
    assign T[125] = 51; assign T[126] = 102; assign T[127] = 204; assign T[128] = 133; assign T[129] = 23; assign T[130] = 46; assign T[131] = 92; assign T[132] = 184; assign T[133] = 109; assign T[134] = 218; assign T[135] = 169; assign T[136] = 79; assign T[137] = 158; assign T[138] = 33; assign T[139] = 66; assign T[140] = 132; assign T[141] = 21; assign T[142] = 42; assign T[143] = 84; assign T[144] = 168; assign T[145] = 77; assign T[146] = 154; assign T[147] = 41; assign T[148] = 82; assign T[149] = 164; 
    assign T[150] = 85; assign T[151] = 170; assign T[152] = 73; assign T[153] = 146; assign T[154] = 57; assign T[155] = 114; assign T[156] = 228; assign T[157] = 213; assign T[158] = 183; assign T[159] = 115; assign T[160] = 230; assign T[161] = 209; assign T[162] = 191; assign T[163] = 99; assign T[164] = 198; assign T[165] = 145; assign T[166] = 63; assign T[167] = 126; assign T[168] = 252; assign T[169] = 229; assign T[170] = 215; assign T[171] = 179; assign T[172] = 123; assign T[173] = 246; assign T[174] = 241; 
    assign T[175] = 255; assign T[176] = 227; assign T[177] = 219; assign T[178] = 171; assign T[179] = 75; assign T[180] = 150; assign T[181] = 49; assign T[182] = 98; assign T[183] = 196; assign T[184] = 149; assign T[185] = 55; assign T[186] = 110; assign T[187] = 220; assign T[188] = 165; assign T[189] = 87; assign T[190] = 174; assign T[191] = 65; assign T[192] = 130; assign T[193] = 25; assign T[194] = 50; assign T[195] = 100; assign T[196] = 200; assign T[197] = 141; assign T[198] = 7; assign T[199] = 14; 
    assign T[200] = 28; assign T[201] = 56; assign T[202] = 112; assign T[203] = 224; assign T[204] = 221; assign T[205] = 167; assign T[206] = 83; assign T[207] = 166; assign T[208] = 81; assign T[209] = 162; assign T[210] = 89; assign T[211] = 178; assign T[212] = 121; assign T[213] = 242; assign T[214] = 249; assign T[215] = 239; assign T[216] = 195; assign T[217] = 155; assign T[218] = 43; assign T[219] = 86; assign T[220] = 172; assign T[221] = 69; assign T[222] = 138; assign T[223] = 9; assign T[224] = 18; 
    assign T[225] = 36; assign T[226] = 72; assign T[227] = 144; assign T[228] = 61; assign T[229] = 122; assign T[230] = 244; assign T[231] = 245; assign T[232] = 247; assign T[233] = 243; assign T[234] = 251; assign T[235] = 235; assign T[236] = 203; assign T[237] = 139; assign T[238] = 11; assign T[239] = 22; assign T[240] = 44; assign T[241] = 88; assign T[242] = 176; assign T[243] = 125; assign T[244] = 250; assign T[245] = 233; assign T[246] = 207; assign T[247] = 131; assign T[248] = 27; assign T[249] = 54; 
    assign T[250] = 108; assign T[251] = 216; assign T[252] = 173; assign T[253] = 71; assign T[254] = 142; assign T[255] = 1; 
    assign alphas = T;

endmodule


