// Copyright (C) 2016 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1
// ALTERA_TIMESTAMP:Tue Oct 25 01:51:03 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
sHZd/YEcmKOMChlevoi/M8sq+BlEMphBVou1JDuggRbGaDdmOLFn5C+xDIOCRGXY
WERlDt9H2F6k7tYlPwgtYsZeSd7kS5y8acSXZ+OcoZ3dl7z+9lMHTZVS0+b0JKLo
knef9Y1E/46NkrUr3tCf1PFKR8AgdSfkSAJazNQr2KI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 15232)
UjpqcLEqinkjuJJaNbFFtmk1nD7z/JCO3iRPaXTEDwFyFjedNA1IIcdOxUANH4xE
rjurqLV6NFPDk4l7swr6TByh1icTS1wEivZg2WminzgCcNoq130Yuf8e2T3dxBAd
qs/O+4IOG94xcgU149UuMZ1FMVotcuipQXiI8h7J3gp/yr6RqEU5ssgvn5M4pzoA
QVd03YpHekF8/OxZBEabrvXSXPSdLmmFPt7AEX9r1zlYA8JHu0hCnINubTj4pKNK
Tzj6VxbryTaIkHeIc5QMiJxZpKNPn71eeac6SV4Z86jIcHh2CRASim+4QCVLF+0d
DIXAvsHQtocczxERTVpvMlLcdw596NmJf/EovAMjJ6kkxpgtI15ZS87M7NNjVUPu
fT3dtQMKB050zR3TXwDUC5rnbTDEPs1MXj8ztk8RoGcjk/2oSZH00dNKTxmlYFQu
iak6dg5+FCDdmjqH++t/QaP2HnIOhJLuxZRX9Y2j+V8rmfK3FQLju0tVyF1smmdp
GR2jluBWw4wyvvzlndDUbd9BRGgHyfqR1RX0mZujp2IHhDRrzNDifCTiHp0pzOH7
rbUgVlT6q149bCWducXSYHXpjiavB9xF/UopjhCCsiblNhnjlYBPEaUocbjgLsrV
remc7F/dhpkCZ/lKbuxSZCJ2Xgo60LiJsT2hn+B/gxZte1QhWhnRQ3bEwa6Q+ej4
D3EjpvY4DeCpvNZLyBhHjZdAUUv/GXPQzPZR2X0Iuugme/3AFOTr6yf9Ct90O/0x
bjnA4yiVkLx0Gv8xLtfKWo5r39WfYlGX+LNvLvYT43gb+41TmoHz3p/sf2lno6Tk
Z+cH9xv0MVs+NMUAIBqL9VAgzh+J4Dhsa1orcKp4VbdR3yTT82AbzxFT4QRhBeuR
HGv6M1APisMBK1dNCK7siOFodOUkrzWzMadxEqLqxzM4LcqyUZatG/5Qhr3PBhQ+
5nNtWPWPNdb2h9zCOHtxDvughDnxGQdOhxe7Z0KYyjbPmRY2lAyCFFG2B+2rGtdl
eZPysiuTMP+qqTIWKrr2gQhII/yqNzntwiSO6OL46ZBBGSk49JPibqMtuwSWmXnW
VyonK2mZxNGpw7MYbvYCjrocWv/rj+wG/A9QZDBEKtCZ2VQJ5g99prmUFe8pVmmT
nlEd14bcbVYb8j5NLfelc6LcyGYTb0spf6K/zuX2zoBImGN7kXrU1xFJwOKCb0Fk
lBz9lQjHjM/KMBx49VhVYIaKJBXtX4d6+mnH7eDej5cChK0hUDIs6zd5f/OhdJtj
tQgY4j/1PbODblYj31evC+jLOVHjOWSLhXj2HDZThgihYx0NldCWAVPkMbITKEyt
HJA9qNaSL3Dhux6YpNcl++3GWhK+zYhzCyzlje63kTfiP3FiE5G2BdA8neJGLzie
W/0jj+25fMgT0btYlpeolaeO14E8yE/Qfw82CckqEj76Tuklv9srMnsk+kBK/KeU
pn3lw9OchN1QyDhuwhpdmTi+vm0RDdmPaTuZjWdnidc27YGeoFFbThWUW7y44ek2
dlWsAk6lrLqbXffjwqpmnzbNRfZkiTQxQc10y3Q8AOYdPdYSYyyuXVp2kxE0CHxh
rmAOtpqFyJLlVLsWgrA1BTB+FvxrK/raCKfTPXXhQpOrXyC6ST18DQ0X2/t0U0of
1jjkS7T/C6+Bgx3HIoeOz3iyACyXtx1xtjBxSMsgzE18IAJfJNn0P35v+A81TMpf
QLocJZC/poskkgi5I+Obfjwqqr4xrZTSKCc56ypY05N7gpmnq5PC7GriT7YgPYps
nRlkk1sSM0oS2ueMB8UsgExSu6JQnQUOUNDU2jQA552OeQHd0KUTXq+RmUJgs1ZC
IJ2EtHvTv3Sk5M06FxyAXhOBPmB5B2HkqurBtYpOsUAVdLhsGo0+aS0x5chgYyVE
atYLGd6uXQ1elON/KjzR8/3RfNcpoRw0FN16j4qym7RxpiwGR4JmSQwU5yxHkl/s
kAH2NASJSN6NKqvTB0mJ/y7VsFNIq197IXrC0e9pyFh99/UqUSppxXQm3VUsmADL
4cLYjoaHm0hFpWEYFQTpcHouqEmM3bc7wWkcgucry3IiuZ3fA/BGmr5K556LBu6P
0hlm2le9cpOe3gAdeubNkoR2YoyNywLbrpECX6XSewplmVwWxxNZiYJhoeEQJRiy
P9FDmToS0038V7F1225RxfyWlIs6yBV4wkmHILDX3r3ybagc8QdnxDD+QfEwnwvh
8qUVz2QlBDEsOyET3WPLpQQ17VZ/7M1I5F/ZvfHQzI8XLq6mffs+CVe7rIkXhZtl
mr6pe23JXiHz3LhpdZye2Vd2IyGrnNZnQoRHYlKj5rqVt08sM4DCk/239ewK9Lq1
alWO3jUGjNYhJETmt84s9MxR42FPDBrk/gMQBsAv8ajBLs+dwRm9cDVIENlwVZai
aXAnZg2Ci3oYFcmUJTjXFrjN4gslAcRVvXrMacjfbaT/1FSMsthEUWZFmca9a/E8
xMUu2iRJ8wx30X3/WN10C0ELWVpD/y5aV8T+RhU+0ZHr3daGk2Dm4kvR46JZbAEO
bKe5s8AAh6zhKMnGit/bJZ1d4nauABoDRS7wapFi5FIVdIB7thfuScUEv7dxClrU
sLGHA4BnQGEett1ivo9T/0P4h5H6uihfxRdY1Acoptv47c3dvbfROeLSHKVLATEL
DMI+B2bDMly45IS1MgIAhsg38baMy4S1hAH8yiuxnkMv3xL83lm4OO+xPyTMyX2D
O7WXcsBl+8ZVnnbtB0okvlwR3Vj/c7ta/lURzxyxdkbGO1NcZvr9qR5gjviz9ge8
9MF+k46Kn4IWgrjKJTRmQHVPv05HdMKUv7SflYK8mA9BiwjaSy1N4zETkpVgcXng
K8iHs8oEibq5k0lYPJsgneujZ13OfPR+bu7vBD9jiK5ngK9UrUL7O754fsp3ZEpB
E22Hr4bKQxqE3upXWeJt3jherVQPvRly6oTZ4Ump7DbWZNGlZ8FaWjwdRV8D/njR
uTexJYKlo6Ie+CYSUBXQiKiYsFblgNBN9ysbPOL5/Jgis2XPqjVOixXNeyRJUbjf
LhmHpoonNOtBdpAEWZBPreOw8z996Z+B7uu9XVgdWl621ypfy5a1mBaXrWJq7Ubm
zzWi89OAI6NtC3eeCBa2MB5Dm27T3oEt3fzahQ6oPJ4CDSUf/q4+Qt4kQFosH20o
l5mvck4HrpsAvqMSoELHZoP2kdV/ZMSMLXc6LunSFnr8P9ziVh31yxbJz0uvSadt
SpSt/gGJS7dl19yV2sD6IWvnz2dncX+1ZOYcY+H+cjHfekhBqubC6UeyDtWy3rfw
Ax+klW6KMMnEIDOST0SJ87aTEBoASIsIUZOM1zAhZitBnug+tFbDY5nFWTCktd+e
4VWI8NiXyHIaWHJd+1KI85ruGwu0dgpL5LABo5hqqCbfl9nvy+4iGY9gZ0ViF57Y
aiFN9TdmZhlbv1Rcqu2jnF1X3kdAGRHUqeBcDt0b70rblikiVcSoBr27eIK3gKGD
dc1/dqBTsqu2cz7Px1+hGt8h58Awyo/+Mnblu8olRIAGTPB2cit3pjzUWzc+xLBV
uGnARy1xi369jhW2aIHTDoDrbiHTqjvC+N6pW++0E5q393lCr0zLMeMZaSzM6lw2
ygFDEH22JXn6YCOiOxV7+1w5O1qrZPj6j4QZjVJcHXAlh5FtfqY43H0wf2av05bW
5ct4coAZjDS45A4vObqybfghXBTj0J36qBGzroUGmVfzhFSGjaVcqvb3rEb2YHcO
eS1qusW+AkUkEJX6c9J3lHJ9lbwgJeldezt+ctul12Tx8fbEfMcJOjyANXy00Vjj
w88mOtjQd3zWSrivlCfaFMlYhMM8nV8rBFIEyeT9ev9hzmzScM376swBDMx+/CW6
JZeNXPIsvEKsa9wHeMSSPnqtR48YLKX0bqfoQIl3vsZvIqZYGOwVPTRyzzDAShTW
4/CwQuVGFu/orHaebVAPk+wf1Je4KdJ9FKrhL0zY/LcyZI+vyTVwBVz60kOJf5c2
EQKcsS7XvPUna6ge3zdZWke9/5JYF3d7sxVWctX/TQW0n3P1ReXwKBNRDca6M77W
8rsryC7oMOvByp0f72h6nQKeID9x/ArrQTpx/OgKYShUteir1lkJmgyggFxq71xK
tg+bXSEjq00lafjX4st+rcw/5vaKmEvl7GMRfHDN+fWvWD1ndEexmPlUdhmH2+n9
nzjL0QqhW3bNiNXMi32QAaW05Qvl9F/ds6VMXUr8438oPMsFiB0HJQJNddVpmgWb
7FJWyJExxfiedWzDGVBsRKvsQS24+Pisaz028s4aNgEH8K05hOy6lowU3+iU+6e4
0VWpWEHOuKUz0kAlFb/5jxth5Z2feO9Pm/iA2M1A4WkmDSVPmkVQwBkau64cGI5k
m6O7brCbeEzItzrNYrbO9xNKvXTCEgCGhXJlQmBaRL1i/K+/CIL2tQ0+CoaEUGUB
DZhOYmRTxjoUQh0zxKMOYftfGA+SKw+ZXWqsRkYeit8T41G/a2N9Wd5Fo4wB9Udn
xIFkwa1qFCmkr3gBnW9UEg/3ld4o0ncVjxdmNAMjis3/ZFr7JIEST+HF7NXdZFuz
TcPvFHVhxCEzQH4s8OXc6NlGyO7unrBT5YSJxKRhPvOluxRtuv7fpoSNSLtEtNhi
CQfFAFQieq7gJ2q2U2wZLlmCKIMyT3bB30aryIbxSZpj0NM9MvqoBhet+E9MFksy
v6jwY9k7W4T8zSqS82rRY7X2aVMO2iJBu8mOfQKxKoA5g1kBjG2QhqKNwIijPNGe
yjsm+XPxo51z5cWoxvONIa1dyQkztur5A0kdV/DW1PDGzNDk53EbLxdQyOFrqnrr
LFul96pYbEku0/m12bGP6fqxO5fo3c8LB5d4+gloBT2fJhyJr20lbbMU9F2XGSLl
rRNXOpgvZ+6obQOzPO6UTA3KGRjnPBg2Enc8VGr/ws+M6ZoZLzEFFwl4EspxA4Yt
Um3OZgCOkbBeUm1VhPEL0R+8k4ah6iUay3vbmbLqS1tUuAEwyuu4CQLDVM0lKW26
DAWiqU+h2Nc+jc5WYHsXTa6lMVMYLgM+7aNX6dQaFcG+Vemkstzj6m8+CUfr94B8
O6klpYDof+XpnL0LLV1qzKzKxfzX3AY9spyMbNtzNFpzdNbu2yzj0h9RRKLMq6YR
3q6tVNUtpQ6OjFiCAKwn9aknIgjx3NdMRH2zNAttuAXcVjbadyfd5kGtu2yDGs7p
3CJsHGN2BX7+Kp7psLHJIEGhBgpTaLs4UW+OWU1lJ+CfdolTro3L/REQmagCo/xv
KBKsgP1FnyLDHRHciDFpYl+JyQrOVOXKkVTVxmqfXnkZXo375QWoJx9IoKx9sYwm
fQHn8j+r5x1wmHxru2V1PMe273OKP8l/5m4V+IVoETFOLwNCZelgdNqK4La2DHA/
zqorFWbt2up+WeIL/BqzXTkQdwfzk5hKBiZAXV5a7W8640wHzUmeeL8kPYc6lsF/
JZMxbEXuW8ZllamiSUURnBwcTXgVKYtQe93Ahrkk09aajk3mCWIyyL1xfRBh/xoO
Hu1qs21t7ogAzItiOEkQMccwFT+beLlFnDJLVWgnMHiqu4M4mMAQG+iNMKZ3NpbG
Lc99pks5DywHXO3/0fdAPRw2xlwSOm0e3DLeBJZk1ZtoCKu5l9KFP6bQSDiI34Ki
CTxoWGczDIiw2oEGSG8DjbrKEL83uwagoygDtnSzk+Eu7mM+BKKus7L1pBHn4+T8
RVpz5/LCVn7blB3RGWYaGebnP6bfBOSzBIFtoD9Xf3yHirAnmLEDgoh8UoKVVWz0
GPM6vx85rQBrx42T7pFr1o9X9k9cSAKaNB/T7uE8ORDDtNNEjDeYuX/dER8T1LuQ
Q/7fuZ/5LR+njGXKkyrJSiWeziPoFSc+xmbWs3GA+41C92XwcI1gOzPAHYyq4YQV
IcuH3E4gzkqlmK8cBiqDlbdhsRyrEUp1rrsa8xyihi60JQiwLeAVI6/+3rGNdjIC
D6wTtx0hztl2yanYYf+Uno3+iIDzc00kpCCHq3z6aCsGvkFuPR4n9wSkxwAs4e13
df7GYFKWINqkrk1fJ1JjhImFQ90eKk2KwZnsy0X9NG3KH7lYDoV2fy3H26jT8Li/
DFBrVEO3o2ZLHhicCPQ84YrJZsGMLSQfLTobDBrASoQNRVj+QjAELXu5TPhfP9C6
yUEAGtDQO7dgmxH2F/TldGoEnNrjUC+9QlxOtR2F6RcAvdJv+7wXXoZHR+KLW9LQ
35yzQ/pLWsMKpeYvZCK/NM8E6tYcRLOHbPiowLoipjhcHU2iRBHGyG89KDN1Rmqp
m8dv5u9qPGmR56+oBQMuuOAu6rfMkGTOH7mG9DYNNixH89leAWiBFAvXhzaI3rXz
JgLPIDMywgztHNeF8a8DtCH3+fKRC1b8wTHyyZh2UHOIQZGpVPZNBFUCA4D8r4hp
5jKY/UXGymxrXmP0NOcoCcye2G9MQFA5+48yKjlgaU98XPPGdU3mNy+cgBf6r4lH
TYTDQvsAm1/tE4AEBDROOspPm8Pu1mmMW3hsf3sKMJsu4Zw2HysTAGXmTT4p95/N
pb1rNkvFpBBCyaNn6pM4LzV43rPkNNIxNuryVprEcZ3eeDbmS072YVpbcaH/L22K
YPkI/aDZXxKPu8w2elVV8nhLWUB3rpM/sds3WJ3jsk/dOd/ik//k+VAFlNqk/Xxk
kNjwcDOBESBfgH6+co4/bcSCA4o2Z2evC7AePdMkyNlyb8ZYvEY2fBsTNlRtjSTH
tAnJrMIzN03LrrJHn0lX5BGiJSQJMNFTXcz60hNQgyznVQmMEjCE7qYJuRlJD0L/
k8VdDvmtbqTTnOIeFCVnTnN7Vc71OuguWd2kHszd+yzRAK3Okj1GcQnGKZVchGoi
ooPDq0n6Fef2vYg5a6WPZYDyk47N3Q1f0mn0kEgdHCKfyZHqcFw39/mkoOWCQERN
NijAucYuyhKbitaYuS37Ck363eHSwG2b2O0lS8wUmHLqZxHIkkAmuBFG38GeXrd8
ExJ8aQiNvuwWW5jnQRwuj897IJ9gkwQNYXzHlZGcrBx/StLke3IHpDFUPOogsre7
G8g3wE9FBBBRoDWzMHoE5RORujPYUNf9Ke8JSwmQhAd4adDu+K0OCBBkvKlc0LXH
D5IAahGnDNCb03HDwUNUSOPory4w2Qdixtocn8g7/gv+0glcQMp6Nq4782WnWL1x
DJWXvpe0hWrwguvweq4AKIHslGdf8n2aAwWVHmQKszIunasufWHvuJ9iq7f6kTZ1
oklRiO0GhRcA6vf9updl2C2vu4o/EKfCqOlY7BJkOGcZQ6/k2VTGDUj4rY8m5B9k
6FUOU1QFO6KYvGo0AIpKzs185bnHSI3jcPcMkQ4+b6a68m0cvWdz60f04kpPx+Y3
f8p75Bv9guO5yqx045gkNlfzCbeCF6WSgQM4y8NF0IdSbsOevmmjj7+68NlHxN8Q
Gt0FiNh6/GuOXTvkW+OVj7V6tIGuBIlXyPmkxEil9/rzWJBcY3FoOl1AGVqnLKAE
p492B7VLqdYerm6tnCNiTrYAr/KNhHnUvhZdBUANdQB5Zjeqrckze+6ltRt7ukX6
AUM7578JLCB1b/3exZ6EXS69pqAIjUXsv6ISuXmIxsf3vBowl0cPDCqQxUH1k2ud
EpjulRwFLzSECO134hMcg0icQFQU8vJXaUUaXnvJj/z9FHFSNL+1qqjaUnpelbgZ
ll7EsvktsiRB5hktYP1q2d4mk0i/qdQGbbryG+CYKa5rPMp4Puf4a/kyBbdCpFoh
XnAUXR0U3T5XkO66fEt0xdLjuA9HgaCl1Ic+kPawHh0Ohg9HgOJ43Rnmvyk0hsYf
z0Ip3Kv0K+kxSojdLSHILOURKuW0pgPFjpSqcQe4l6axk+Mg7v17wrXP+Fof+F5y
vjH+9BMf02zHiPa18x5VYAhRrvuk4MS6p+jddcVuOc32wK8g+h9CjyB3GH4/HAsy
8haWrUJiQVvi3REE7c5ieQcFVOtqJay70apggCHNQHME7nP4B85MOnB9b4NlXmJx
CABJlIfHLhXCe9sOw5vEJV44tAYMPpAKucFrWd+w5KHRWKjnR0kd9owMIZ77MxTt
fUmAz6soFDWIdK61BoEczhJcuk2wdm1h0gC8nadBpI0ZrQfL+cqEbzf+KUP3bKc/
z6S6WwO9HEtcTCsdyx4Wbn7/235wKYuoDxCjnH/mNpnFdLGDbrU7lJC2nlTu9iBa
JUdjJWA9uV0vG4Zqc65yRwcKkUZc+TqwkH6WrLQKx66EDVR9GdlgJz9ZNcTTP+x5
3wZT88LHY9EbeZTKdPzxkREUSZoANDhbpEFlMziQBzQwuFqwn6EPrvFLSYKFCeKn
xhYqKtHwEhbYkIhyNuzMXNaLpYzmK1rt53ZrPBXxbXt+wwxuL/Zm/pK4o79TO9Lo
7lEnbMdBtc4SIFUgk3BeZAmNUrESK8X6+osw3wIFntoHeB6h6MGK7HzuHask4l0q
0/ySUZFQ/KEQxqSoXiN+7XSjRn0NXR7FXOML9sZQBLy4b0oSVxEIbQ+iZn9U8S1n
A27vII1RbFCLjPYUC0VBZJUhXxPlhGd7YXlOaF7HyDjb4FBQs8yCgmnHYHA4XKkb
HnN/mt4Zk/U16WWWcpnyhxte2hzzLRRADNhg/0Ox3ItYJTPt7jZDdXa0mq0sX2Yw
+h3oB3c6zp5FHLVMnum9/vvsozSdgAjKMIP11bFYhRKLqKJuxPgNyCL50fDQTlWK
FSnBZ89zyV7NcYpwSE70xi69z9TRYIUMN2qwWZFbMMif+l0EgoQDLtsR1Y/7GQOF
XsCvLhigM6zcvBtdNxPT33aeKgn+tYK4D9Say3K4NRUpQunOfj+4A83Y1HZ+MjWo
ZVJpDoHItSiqMm2gXnXyIOcQQaR5RSKofa7BnVElB04VQoyvhKS9zGrzGEn2WjP4
kNzBtsC9UAHB3Oqd1H85yHjBDLygj1uhQSjGUCvnDHQSkgnIew254voDeajnOw2U
KK/7zP7y6auFbHbqHDHKj0ULLNyun2CKS8E3vyZKplLEzIqOHMQqXwI0/ecbtyWy
8eA7YS73RrFzDhLbBiMWIJtS6XnFueuE8QXZXEGCy2G8cQcIZnfyjjZi6nY/fn9U
ur4pzn6wn2pk0n6QJY3QbjFoeiCBeux+WR9yAYSbVm7lNlbOV281eTCQWLKBBYYM
ZUzkNZSdWsvnN2qvazOtUckDvfs8WdNzt+XOQdT4eowT2Qz/l4Q/HY81hdct8aPr
gqxqBaxfPrA3zAGltm4KSL0xeARL8C9aMznkAgTerKWnAiACfgPqs5UJP211Sqdx
g4oD0wdjMdwiXfHhDiVO9KsJ4riu01IaEtiUmQjH0WFWbYKMijL1gpC1J2Z92QiM
BmCCiXr+HDYPomrt6Gfeyw6uRcRHYP90pVu60eifycm0DltH0LnAklCLFEVfLJeH
ZcyA7rVETCEqFXePjunaT2JIozzS5fBWtswIqFAu/UmLBRuIY47adyyDdRddZ7FS
v49A8r9HH/JSAHIWwyyZgNgEqftZIB/Fr0TALhtP87Y+Q+qpI9CTOgi+6Gfyl/bS
ycIyhRGcy2XWrjSWMT8DhoAoagzLWN4D0isd1uq/eWmwUzE5gS+5BnQwhW9oBPyb
EEqLP9+7p1DGLF0qto/lhWtSGbRh5kl4T6ugB7Isb3OyDhMYKwLuLFXK1jZS3IaK
9VVz816KLJ0H3/kM3dvKLXWa4L9dKyDV/DeTR3g1CGATqkjpQf7NfVJc8V/9L2Ug
Um5agNHbphHSfP/jqWzVgo/hJv/fTMGGV34Qgo41dKiwcWEVuccUpAAmUPjaw9dF
NmIZ+c6FjA2e/GJ/xA32mCECYRftQ819iBsk1428SM92uQvYsVGkbxmWoQdhHPEH
kxrcNyUAuxnNtgYhTHAvPHq7fCIhJA3nvrrZlPFk7u7bjrubk0nKsad/gnmNqQrg
A6vN/qOPCIb/rg9iH4VJzNqGeI/HU4u7SqQS7qWcRCRDCCYo9DPdmZufQK5RBg6l
L8BydqgZwTNspgaI8JXYKLHIHVcbzkTc4DVNkCYSXJyaecL2riBBAzOhDzQYKbG7
br6ixpq2EqxAYODXlitY+3vth3IQgt6rG2A5UFPYJNGtbyTh8W83xVKBeVZEx+1s
/vSY/K+Uya9T4PcH1yeCuSVz62bcS3TYtiCJ7BWPADE6bnEusg9cI7zvnDwgvWjM
1Re5M7zwS/6ldvk5ShTfeJXt6z6gf65hEaT+XdUDvdrhgVHWNkYW2GsfcX9p64ic
emNujZjGNi393UufGIzPoZuovzPpNJmxkQvpjcRHt8hdOME110bg5Oghl5d+LOHH
3PQc+KFrgTUfRxaseeaR25m1ubR60mQs1FxdLQz1tvQR12D1c0vygIeLsKGIgjsJ
mddYEtVEM3uhMa9jaJugnp8k4Xhpo2XVqKOx0U+YiNVCxNMmn5CSTuCGoS3qQiMn
IKNFyZSa5JF2oOeImw3h2KXUjOzOACKymrMLGJT447naJR626T8vulSLFLTh3pj6
W6rl3m3LXXCL46hXNpIWcNXzpzyN7xVwD+nAXLn+FPd1DRA9i3dj3lGgYPfjFhYL
joiWPptD0dHVJPyzjXDDuGa+35eURJBg1kDfX3QxQWbUEwiovicue8c2wGpjTH92
B+dAi14TXnXQlNyh7vgsss+4AZ+0Y78FXUuahIuNfYTsdQgShzmNxK6v2Kluwdf7
A0b+wk7oINeyJe9yk7j9tEO6AiXI+OqA2Sw55OzIKR1M8XleCFqm8Dl9DdA308S7
GT4wCDE0Ey8tZPoiKLOfrNtOPwP399IqQrBAgDdNc0ZnqtsBwNfDpO/8W3OHlf31
Id9pd9j2+xBgKoAtbt6M77aHfEiBEYT7xOfSJplkizphPax8inoxyZliuTfQ87Ls
OaobkL5zPWgmw+vv4NXafdQdEh/GnNzEHhWOlnUOwzmk9OMU5EutmO7EDSFzliO0
mWuiyTpzbrSzUNf3Q4SXoTGtI8iDGA+5eb3r54NT7S9BfnuzQ50Hj14rzgJwlVpB
r7noQ+c1i6jRUA1eD3UJ86gm2vkXQhmgPGDrzlooiGo+QszrBOBTCxwOsWKnj4Jm
QGP9edM8I9Icmh5Et1OuXLwgg9Flw6FgCMGbAZhrNwDZM2JdIPWNNDmixAsN62Gg
aMJe27bRkBjoeo4mvxIvX87b4hjXmEEN+bh2wG7X6SIRNyuEOj+IFvLxT6nHVnRq
e1+V073mdlPm8BnH5U/dxhpwLWN63mJzbXxKnp7FkIKTxZZozCoc7LOHOqy+aAyu
mwz/cB75wxnlLEVHAU2Kg6U6CC6n8vRz0EyWKdFWewB72dIRzMUFB0wVdmIL3HQg
ePOgqyr6uPPiT+56BgnThsmugKl7yjRH4rdtBbfNzZqR9Qlp+ZJ+VW8sBA7IN93B
ImrIAa5NVceRIhYQojM2I4fGSUaSHPK9/inZ+B5xq6Ez2gB70BPU8FF6e6xOP8R2
GbRBliipuZB9Nvq2vpOxT4afAeblCEiJDpHvzQPSqrUgctQ23r6L1BD6MrI0kRke
rPC4m6vffsJSYnCqrZrneqZQgDRJZpivhbzmQvIceQh58I4vb+224D3wCQvUBqj6
+i3KWf0ncnh4f69vFW3q/4/Y5yhzksZuwDtUl6QGULvJQkHnnf4BPOTa4+eS/3ll
+Vipv4kWbW137bbhyeYQj6swkVlRuPczHCX1T0uGaN0+M/RYz2hLrnwwwZCZlZjU
IEtsk8eT16SmL77GYhrQ63At063ZrrnFU5y0MNJUwNcnHTqGS6xyhzI4BDE/AtOg
3Qs5SIMVEJQKZ6/RX+ricYAazRZSWL/7Zwzy2CoM14WK3eq4iYLa97gG5FtSCXA7
KOAsoLLiVHWvq8D1w6BrhXSoP6NCKRfahtTfU14bV5VO0GMXy3H6+qoa7JP7CTsi
KsxMaSGYSJGgUYiA3woA9gr4uFUlFAyTpjhQb/PDd3VJvEC3OhU1kNnUqKSYTZcS
gQ7lZHno0qbN70RlehlxlnJjw8cW6npNl05foPsZOu9KEJXtruwv8SifUdJHVZfV
CllS2DveUrI3pyq+JNplVmdy1fa4xTVD6ca/AAqRTd629zyb7DcruaTkSvnmzgHi
4URffOTufkihkgNRIz+aROjlDcIz6AW4DSTaHRd1sGGaNAPKwkWHsQ7nU7MhqEgM
JX4DVNZzCA5uxr4Z71n0TKYv9Hd7NGxDi8hG2o2YvT06D+bsTYIaJXLVt261DK6k
MJX43+JKsncc04Rw4WsEga3ZJcp1M/HRdP9+9yMGJ9FigEXl5pQgQMjjcO5A4k+V
JJ/HY1hQ5Ee8U528LHbeKxGz1JnTPVN8bPixv/917rgPC+RIk3BlhE9WFcsCsIxF
SCjL6JgILu7XOn74aD+5mLCKD+Gezptb/NC3L0z5Oj7bLOUcE50C+2qb5nd3MuUA
OyLOfd2rOpoExPiMoxifFN4ivNL+hL+3kytm/DQXmHct1Wt4Lvx85RXD6Pd7dAQ8
nTdcvoj3UgP+SPlSA7r/Y2tKzTKB80MSrwbi+TOzdcDXaS7uvmdIzauyWPRt/Fi7
a3I62j+SNaK/Arew4rhLoK8habEJ2bqZ2Yj4YewSrQygPZlOEHuIdxzQfdJAvmXI
X3gIhPZxnNJv9M7l/IU9qyL9JJ++1njMibCzIJBHvidaST8ZN1WU1GDPTwLX5HVm
JWa9jhxOOHkUalUoUKEubiqk6iUJIMMPmA4TXGTqPtN+FKWuucP+wIYuX07dJdgL
awXEc/ePCN9k4fjynYmZtwWKtTyRU/760dUgogGybpFC6Q3AAgZi9jKEN9wwsmeK
zx5x/xPyYtF4WQ/IE3Kq3rQK8CofbkVW9rLDNRC6I5hQJ7XshE3sO5/0cXUXtzCM
rHK5S9AlZYFRuSTFqigGphINi3JBCS8ilYvXh0Pywx/lOsCBrL/rI4syqRQ0s+Kb
4NSfrzwJ8onYxK8qSVxcPnLmmBTQmgPMO6y9KE+BDXNbdTRv1KkOluEoCsDzjsbs
ru3XeRGLRDvx3nOCCiJPY9K7b7cn4Glhf3axcjrzqWZVmKsHkCzDACIUlBbJYN93
mEkagipNN5uV3Rt1NV7jR7x3fPtyGfWmPVX1HwqbG3z0pmCs2v/XyRPdlICKJolG
U0gMcg5400vQDa7xtk2K82uI9TZOGY6H3e67kNALdBVjLbYnVVy+83qaugzN8X78
8xNqeBo4UJiUCrXraTa6zR5PCrEWFaFkkAAPcDdMKSEQi6Ge2aS3HXQaNLb6ufgK
723GPZwbh+A1yWpvcu9t5dmcfV2Em9DINh+7mFWSaSZcPVdjkS2ea5NnjXrq6VQE
w9dEoxW4jtk9mHfOTbHeYOFP3Yt9N3XBiuxKrOQY9ey+6hvA0GTdW+V++Fhdz9+V
3EFaFUxrnhLujs1zmM1L0swQwP7JXaBAU0OcEphJGt0suXuUD9zGCmRFaTWGI45Q
yPFL7jvvz+NFcBVpEBHtq2+ENa/cSjUig+EbnvGEX7tE+41X3zpsdUyOlpU5ikfq
8AYQKjrBoA3PIX1cRQnj+gKwsWtYaawq25+bdu2iCQZmTzdXktp5l53HrxhaHyRp
kJ6xrM7LjxMLraucn2w5JX67DYANDNt7RokBPMZQKxhD7Ma+xlsouGjlakUo/9Rt
CbfJR0cd4vj1LF4Xdsd1k86n13PtoeNjAWm0WVfjFW/xrhRdZCaOkJPentUSISqQ
rc6p0n93bV0nWIQWgdkWa8qL+151F2j8wazYrLu/c7k12Cp6J/o8yhhxNsYKkQ90
RBHxK+oKl5VJILcUCGG9Z4A8v+kMekNAjoxEMT4b6uzpR9b5o6KsIWF+/Qmka5lZ
ao1pyJ33goy1uCFBNZPDA4qRXmviI8Ctkr6PC68Q4VkaCgGAIccz6WwaawD37xC4
e91IF30MO7MAkRWIIcLeZ+ZrmTvQfnh5NCDFXoTbdBT4ESFQKH02+gh8YRYJb65j
rQtlrc1O/0e8RFVCzf3OGLDc2ZJ2sqN0oeJIpHDPDyHrMtgbEQV1VS3uQZIIgYwG
2MuqS861I2chA8HO9eGmdVJb5AOUC/yAA12S8fY+IgKZMHBtDcE/LUkGxESHRu1e
cbuzswczf+ypWeFn3Eh0i+akFuKvg9Jb1tTGyQc/4qMSwy4nVaOlVHJTtM6dBD50
3CPGo3ltnJ3s54fRZArqtO1+V3WjKIdiqa/G6kD1KeTHRpieEDUnMwy1R2dZJPUQ
dq3nfoKPAYQ7jJ2C5UipqeL43QGmdcvMjGnJ6QA/VIfNkQUUNFHY2IxUJKmVdQbo
0qz3gI6h9M8ctzODBnS6sEdFazawk1OlrENxytDxtcf8bBDk3DCckCYNPS/FNfQh
4cNuO7ngNOokK0ezrnSsLCvkQ84cbY5bsH/3kSRFWNzrxZXJqw89F8GWij9dY5u1
EP6Iu6CIe4/H4h9HcWPaGO3PRm8JLvmwh5GQvnpLcPNvBHVampB4nutYbHaSd72V
sJGCUZYKhMrnIcl8ZH/zOS+NcXTQADeAd++4T0CT0jBu7Z/A6pq+jeVmAS6BjvPm
2bmocAiL95v2ZD2Cx71+iZFuPAQ2zX+aV5mB6n3JKZ4sajhjhEqvrdnx180yNOZy
seGRa3H+3Iv5dLjKdqY6g4S7VuieBeDTgG5wc+y83e0JUGeMhIIact2aD60M8t9m
mLEZhLWaj/Aevw6xIlZUk5EERWSvj548Q477dJZPLLzGArhRkrRULZQhjWUs44RD
WhO0GH+jBPIGOPva0T9OBmmlwX6IopbgL3vbTGpIpyDdqoAjGsNEGpyIsjAc5GB9
z6g1nnPQ/gsme6zCKB5JqTD81/jSQazTEMmDOlpTrrtneoh1LuKnomvl2CRhe4GK
g7aGYizuK4i9eZpswosOnxO9ZmiSCEZ6unlyFCOdDLOiwZqvQNVoU1g3zNw47wFS
uBBnYwOeEV2AUwkC+AsPsEyVnSn67KJvxCmHrssGI0J+UZxvtFwy7TcEeOyeQiqo
MdYGHeaWGdQyFsDsBObeIxq1bJIAG4z1zR/jABRWesLatL1ffOK0jAKYwgmaki15
9kN37ye7+3PQVOnrHadbZk44yLyJQebCm/XXCPrsqT9a0PFTLg0O9f06yu6eaWWA
OHBQJRdKMq6bCfqF5eqxuEPzoGU8Fo4FsQ8OlB/okmr9qbp6U6ZpsrsnwMHOwQI3
aX5qqHghPX32kWGVJwQ25+OyR6SWl0Fhpfr6s/Y2iMqx7uyccqp33vxoB8luN+cQ
Y4szxC1U7EitZ92liq80NB43GNz6xySGIZgHYlHuldwGu3XfKRWxkW+O/tvoSiA0
ATQKv/iILGXO+HeNAcYT/I4EUSjG/LkRNVS2VK79xOdclohJsVmSt4Z5U3Z6BcUj
1XIMmteQZ9PdvOua/VcVBf+iCkvK0tCIrFt0JXWeyaX9wlLipB+FKLWobgOsQwpJ
UAJk9Si3jvjltDk5+GQresY7pU81cNeBSAjyGXLlGoFVhK2etVCM70iWaGjoFkeZ
aVNbOhpeYepFEwvGQ5T1X3DeVlCQyfsH3qwRxtsTxSgBn+LxWvPBNqxcSSiugnq4
8sGZc3ltZkbOBxY977ckjns3Cw6WoMsck4qZWZQISGMjI2zHLYtzZT8qsp1Zla6D
cvKzmg6K4lbohZKiPcJhfR9hCw/1TgNr0zb/4Z09gQLehxF1Z6t7R9OhNfGuKUxF
XJUbX2TQ6+B2S84Ul1YX0NQ6KNqVoBZOupRrDVJjwQl2KZqQmi8ehWPaRgE++SCe
nTvxQ0Ug84QAK+CUVJwJLJli+omhWrcM6IMn+IwXXMXl6c87m4DQ13Tw+AaYftPp
y+NVlbM7nLZYEEdBwAFxHlPTvvwKx4/9q4y2vjPcinG5ufwZxrbLQgEs7faUo7mq
80x1+pJffX+2PiB11lmgmKIVgtXoBc9r1lLd5OuCn+dZvHpL1Lci+gDQ+h36X9vE
Ft9qFiDQnrYW97CxzwtpgmPIJQ4uWQ8TlgjlPbnw2mQ2X8Wc+OJtc0J/wGWWf2HB
1q8fA3FNfXM9sV20oNObBeNbq7n7by2Tln/d8maoGR6EZ+SAbrtULGIthm1XspF0
TeM6JEqOj5pPZMH7eNKWB8oH2e/2Hw2EujWyHXA6/VrTcqMk4k2Y1QyUUFuEN7+9
2jHbhn3FrBMtSI1lv2KieoeTqe1OtEIZbuy69RE8EpfvMpdovSqk38Qwl5xe7qpr
TfIegYapNpnRdfWWOOCqL+FrAnTjBaT2O6W8JnnMzaWX28tujBMcAqeSuvWmcUYL
uwOaK8RkxVNZCG9c1CzvEWQ0bFe93FqoH/8sp/L57cA7qFjElllo2szH4TYnTU+l
HrDLe59bQBkY21cxk5IosLo/MrK2+tKvb4rlXuoBm/y4xm6kotVKIQmVeOYZqZfL
sl/1PmKr3g/Shi62ii8KYBqb3A63BlMzxkatXWD+OKiQMLVF4g/xxx2ynLwD0ExH
rqAZo0FkjYVI8GpRyTQ8uMquj/JgexpnHQwBhdZTCNI4VAgj/2B4w/JGNuWeIJLY
f2a5o19ZyETB2HFeYEVchwzmY88nh7wzomEFCRtBg5pQ8NFzXQNg/iUlZ2hwOKkv
2Hiniz90+3GoCg2FqEF0d52pvENA/NeNdXNINaOUA5qpiqJ7KkVsHaqhROq7MrS8
8shjHI69QSsDgsdW8laolzQlT14SBCi1eyJYZwkSubU7iYvJt4qWb+an0yyn7bJM
82NtY8M3H5jdbe9r7lZNrHy3BeuRFiLtQNF8Mg2ySMk3ESQXUBt7iYXU/60vKpFM
pz/vs15M2i/Uf1ScQlJVkrUR/MC5sQTrtEy3XDBfvCFDGhUKf+1gbtNgKSRSCEFP
jK3jYRYYqkYJ1/yC2TmQYE78+/riGjEzbGA2aiclFoMNy5yxqZWcQSVdYMeIA+2e
KwEzQ2yhAsiAvpSlgkWqzIWgEwFgxdijc3zIMoCaZeGo0pEfrqfjgrXnTlgCT24B
O6xI+RUyR4jlwK7ubJHj+FUjNmJ1KDPMbKV+nu2oVXeisaMqVy2myK5BvZueV5Of
JWwUYEedQWyWLA/0aXnt9bO6rNufdXL+8lvtsrMduRHFrqj/4yREU/pIeCPR0Ovk
B5JJ+qdbOoyjVD86NMFljqrl/yt8eeyirXH/J4ul4UAqFXltvUddE48zemdWCP1b
2Yx3e/tXbT+OO0LwLMOPPMdUQA+PxPVqR0Hd9e+DtxQHzNaT0vX1o8Jaor7T8LcE
YC5kFJoe4jGbzOg3XkAeJ/U6yen9LIZiImNpphMEmLjV2/ca1WJmkEf/F65DlGOG
5gWcLAn6VtVQ5jDIsIB2WYDN2sxp6Q0jR0xJE+tKZrZBXHMFLLVqXVPBcX/121Ac
vEiIivHg+cdxP835B8pj2QL0rRTQe4VKejKJIoKOcZmOL1G4LvI/CIS8QJKdYyg3
jUdwWIYuudiB5QPRYe2HgyfmQHmEEXBsNDmXFKP8bSubhQie42gvU5XQky8aDmyY
rEPFyUQZxiBIBjPVbew0Apv3EZpgIw7op2AOvdRsLczowAWywW3IEt7liFgzMKE3
zMpMdI89fVRe8GtNdcTmcc2Lzg1LkGemQYYC24seQDk6bUf+eAvokca14RzjnhHm
lL5/2nZtHsLxlhEEe9LSzOV2j0uzbbg4+9GL3lRQMgI5EAgEPOTBmpK3qCiXs8a7
RRR6peNWjlTrtuRCfdayyWIFdP0TzrqZWicF7JwgvsmDXlFZAoQFCd1hmlDr/n4/
X8FqBiVanIZM/dMf+uIPGMdXM7T0ChmWxca5LhKfWEaruU91WwAI8TOZYxduBJ7s
5bU5w4cf5sKI5vcgh78xhe7uQX4RFn3H5F3K/SOVLg3GmhfYhgvxsrZEo/RmsYtJ
Wpnz1WNuEg8QV57fIlCYpQiNqxrcuL4QxJXhmm1zFjPbxGMjBBNg1u62yKL8esI/
d4zRAi3Rm2e/BO5HGOnSCxprwDk+0kBIOM+bhyaJ/dqkUy2Zj41XEx2oBsvn/5fC
R01mpnxHzX/h4w9iKm1QZ6OdhS2hNzxmpcEWt/zHRNYmrlez3WURFJDpR7nq3Dkc
15jGOerft8qkEo3vWuEBc1XmIQLd6jMS0y+XWX44ZUejGIdElRmWYM1D7pX7s4XW
Kmya784kIIg/FBCFx/sfezJtpXHwF+HapdW9X6hCbiyzr6lO3yzac27e3X2+0gjE
lUIulhrhPFnqJti6Rlhhlj+vYDgY7ML3Y0TVeOi4EMN1IbTKZmudtL1cw0Us3kZe
JxZSq12FcloA3t32KwkWmtN94dQS+tIR6z/X8Qates2Da4eFbtxZfgh6IzDtgnUs
aJHHvF/7+YgFyvIll0wSpYXduJNxrYdPzGLmExvMMxGdUiI8dp3SJpCDGj4qYyAO
TxW9NPif1H+YVbUteGtKbw6ii0q3SChS+l3XrGYIbbhJ0CkuaqG8cGax4it+NYLS
+5uAXpuhsgjtWxM7cSCH+rrjKsvlGR7vJj9kSOodVI5HCWOlJ+ZpzgG/zB5DhnNU
WwwobVHIdqr2G+WCsgAjvJ5w6oDDSpqngUTEsj7Lv/T8Eem0oKXuJmE9PKAfjvrn
jFIrHPSOF5QlgAzU+XxWFE7V2FCRLIMlJ6vWuNgJuZ8O6GhXI3bENCMTHCoPd+S6
68YAApBUOmdYTWgm8qn+HjNqFtxEzkmLFAN4kSPGWAQ69hg42dM53pv1Y0DuLxce
2QRbboRShjcz4VQFIOAFUQkft8gCPBz2FUCA1EVOe498DIVnwJw+OsrunglGXNtI
RDdshZdTO6hlDSdPwYYEnBVP/sAZJoeTUd+tOBKdnqa7WJp5JNZ2OdF3L9kGDTdp
aE/8/VNwX58dJ+JoSlPeI5MXpuCRa4Tsukm3OP5hQCPxJesx2szmsKlMW5rELN4o
856vR7Oa9K0Vq/HxgTGRVTa7ky6aDDMmdcjGek2Lpt1BvDKuvDaZq6YbK7VGbVzX
e4zjlCK5TqE3d8upqH+n2N1TQ0w0MzciH6skZFipD5+BJLkluOsLU5vCz4x6hLU7
gC5KuLVhViOTCjWy+GOrYuiYbalxbLzdrYUgWOufPzcRiEaz5jS/iFkq+Dhag8/7
n+0yw8kKClBCvJ0lnaSSaatjzDWZ96hMqUoXzYBrmE/ko/OCi0OEUESVd+GGkNY+
lllyuH5EFytJTKLXreFKSutbmrKvDFCOix0EAsvgCuvzJZfHpNikCu9SUwpBAgyr
n0WJOdP6pnIzKcnul5sM1lCo1tG1x02wxoZdJBcTZojXsAzLpmhdL3Fsw2yzFhVU
DYtaR/mgvrh/yptnExio3mddWG+0SruksPwp7JJOjsBbBrzJa7d4w6DpXheeWL1m
PN4Np5JPr2JkZnDSwIB91vunmosAtRZ0UmWbvZCLO48O//Bq2YpE704owAldsrBV
pXO4dtKbW+K3Z+d9THOCgr8yHcAi0qkcE8Jrx90V4XmdtFerxF9u5v+rNFdfJkiD
HyQAFR38Ej4FlQQv0H+Q3fNXKWJVy4D7EltpxjM3H4YsK3H+VUkZDzwPzRKJIy6h
T/XUA/YVd6iR37dkyBD9gwKUMhbowEexQZe6pSQnPac3jByIl63bC48kf646bwii
MdRFXVU7p11ERaOOLNi5CqyPIm77FiLh0FysYSO6R9s9cTBbuAnkHxH2ixxrAKug
wumqXJA2+Uadxq3qIxFQg2f0c2ex72ImOQsDMK0NR5PUCl/PUXPaS6Vs1P+zPtOq
BBK7Lqn08JN/fg2dk8zDbCpYq+nBuG4sCWWHMir2qNx8Y5BtptnmkxWdEU5fB2aC
A4XdU9w5JxaIaazzdXGjgssoM7nvcaZmCQOBL4FF5Zn43KA9SV4V6I9wvaS0YvLx
L7VdoloCMJ6rfGMaqil94VZ6lL2fAYc2aXYen3AcBi584aIpof57L/FKAxKSytA3
QV47MZ/hS+IEB1DZAFyYuix962nEnCsLrbVKuRl0PKp/5qkkErxtOGBNYkVtGJ3Z
FQq3r2lEtpPjud3uYfvwl7DQ2D3FYlcEzIdKSMA4mXP2ofuLzhx8bj8nUumA9FTH
3WDQmgnHSnM24L7dN1NRt0m/k1AM8SCtrD4CVW/I7JJaMMflTi2nPliPTu+OkBkQ
ZEr0mFeu3u44aiSGJLqzOWhTvgxQIvivIJghWbRE0smEhMxfxNnNxHAMET4AIJbW
TgEtjGWwPil+K1UIYdNTnekGC7nwLP5u6udSxyfGo4nublmBnyTJLx3k9/HMxTLJ
u9Q7Z0c7xRoodgiSLqHNRQ==
`pragma protect end_protected
