-- (C) 2001-2016 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
F3vu2YmK0zOPCrw1X+d0wWDAldtrVMbpn6IBhoaSo16F+jTe10M8uflGKJCJlTebJfJ9E/RO2eX+
5XnQluhw6bg3S+RZwyE2TjL5g8kBtErEFY6jCneBXMbTGyjHKjFjeYtELys/SJZEyjvO9jQB3yyR
VJsncloZy3ctj7Z7pLCMEbFX624/8z0Y22SLGtIztJbB779B4DiVniSrzJPHsK7p/rbGNJdyvBMS
1oB4Ln4kE7XjB2UMRoK/3KdJCVZg3+zmkgL/RXiaYe9GK27W5OhsD7CAHQI991lmtbUdGDzMWyG8
TdK/qkBVeVWFMIpe2N7LJWdulgObZ5bGvqgB+Q==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 12752)
`protect data_block
eDDLad1HQGL4I4iTrOwwTQq6clSaLqu7GPpReYD18WtHPWk3l4WNaR/sAHWzv1snzGVk4Kiy0yRk
zeb3t7/5cW0G1qh8WhM34HEa6wNB4xmXRH2xbUCTbri8VJjF5Krk6/iqZky/gcxor3xI749YHOrv
Ma7ohbPO5y+DrKv1jCZVvDZKSX36GHsUF5cpr4AhDzoORHsWnVtb2HcxSu7qG8vhvhx9GRFntZYx
e+zyb5pkaX5bAn8stbp1hIlBq23Np001XoF7PLBjUbfh+u21IwwVl4xyObm/fs98QR2cU/I/49kA
joXX7vBe9uoz2ROcB0UUXKzHaZVDbEjUGLQDPqaLW7Y6XlvEVlIh+i9tZIqjxWzP+r/gBKcww6Im
/O2k85OBZUgP/SPx3SkTSH0mcFc9aKfO8vQ6dO9umuw2vHlPl4rJ09uEkJ21pQHl7+ZPXO0FQpyl
G93O8ytgX2GSN1AJVlXI31985vWPUW8YKhEqSRCCe2h4ZpjLobtgFHeUmvfa66HXNwGyaGYkrt1d
cl0hbNKt3k0wV/tPDF/57V0bYYUbamYYd3FvMhYABK50EUK1n1uZRH327Y9CHGpAPKLCEB8ut6lL
6js1lzsyw2igRkpkvVIcfvFliOyQteWwidxNCEeeQanSE02swqvcF6ER+/A/Ov1/jpjFiSx8mVrJ
x9TmbRWjk7zW1cL/K+4FuWHpQ3b8Y2Btvj2gY8guolWLEH8OD+SZSEX4QY5s2mPO63xY76KTlhtH
IZYwFAsHICfi9uZB6KhyDQvRK5MfR/SD/E6lh4ig+jXyYk70PiKUUC70zRHegeR1FzJr7k1nsM9X
v/ot2CfW9qkjbuYEv+15CknsjomA4ycdUgCebd4C+GlcNHMdCBi0wAfo1/rBiVA2kNBlMcCbW+xS
QQikv66LrJde2vNE2i8pBI16IMR5gRzXMmv2xruEhGCGXaIXWZxl/M5N5KX4Jq9pKRjt9IF/Xhq0
bsjzNOG1ZsgEY0dpal/yQx6CXOfZozgygTgkyyuKj87rCNRr4T92KZB/cMt5jR/WietsaVh5+Wnb
9qr126NKTsRaV8YfNbgOb2xNhTF5Javfb3LguWkJNG+fiAU/3pkb5TZq4p2aYMJf1zs+tuxtrY86
MEJnBRNkasyYNNP0Eq+RhFyD9zgXZvh/wC+0EdbD16vHbaGEGZZ0GcA34ZOugd2MvjCc+0lIq4fc
1KzPpaAyfF5y4+Cb/5SdphS5Y94m8pCTQRkPaAU2ZoMDAqCyCQ3Glse2tPQomXrltSpm9tbBNihi
3QpwjyyuR+8pdeidRr43qKPwYAFP/i6ZKX0MLHjRmMiI7Vlgh8D1ub6Aa5tXf4ZHDqSiLULwb9Ck
dpMwkXgjY0u50yQ7kz6/0TGb70K1Nb79iHcTCNDoxyj5YdAsvP7V6YW8CzKNcpGY5qeoeY59NjMA
dXISxBMikjLOefsSGf+0w8pFjZKPELpfPZd0rN/XqmBIKLXvXt+3hUmsp4y5JHKqZ4CrCjfhmxqO
mZkUKrt0U4FrVsDc3UVPqKfx0iQv4SWavPrOzIaPj56YVLTfm5v+Bxa4o7eIcV1SymMpLRbtj4UQ
G//xhSpOViNfIdH00L0dhZf4kZZPsPV55L3fIgVOWghJHveZuafbdy2nNrNz3bDUwKg+9U2H2grx
xzomKxlzrIgR3S139pHMWxDOuNLM35mZaj5gYWb3i3vJN8v4dKUwF+RiZkuF2zZE072L/c6ZWrqM
alTmxtkzB33asleFrNRHD6nX7FDuBW5kpvHPL242L3kPlQEEdYrtYbh1yI2j0ZY9uzxuTZGvygsa
BD3BQQ71TrBS0hs9Z07gp2LL5TiVgQ6jogCrdHk6QN7rYfXioGCWojqR1y2iYy6uXqP50kKxmVIm
NS0DAYLTFaDZGCFh45CVtxNh0xZNhFAHVotlssplQX2KCH7YGjVIOoaFLUOSP3I8Wfb/mrL28zM4
jlfRvxYPw2ArhrM5vlWnKWJJeDwjye0Xa2qmMyFEpMQJTrt0C2v7way9h1ZSUUzRxu7PSGkPdRQJ
W6ldZSqd3T/VZcDQyN2frtCyHKdcg4KYGO8SmpTr1LjnTH1C1cMMf/vYrQORCnki4LZMcV3jBkYi
XYVFl4gmfiAzY7Ve+ayUtTFWTDXxdaY34Jr6CiW59KfMqBHrKNz3zw2tkIN/gyrJi9/OEQswFDPl
39oIdlOH/JTOlFNn21OJpX1+rpU+PE5nXRL0950lOoxvLfxIfTOVws4MNEmGl8goNyPnrEx46rn/
eKD0kkYg6Ag01y+tffD9H+/dkUu3b6pg6J2MYqWl10/urWS8v4zP64lYNxLndwfJxtj1FtYL/aXi
JLHEwXDBtYizOZIzJx8QlxyWRUIgEED5vja6goeDGPffTxI+5j6mHyuqioQUqpE/fjlQQhW76W3i
uQlZ45qkEkHDBapRkXIlYJufwnfJ1WQGYZrq75fmwDVDJjLVdZJmVF8yY0qNZkBn6orcxXEEPe8t
WmYyAecjL9jqkYiyzEyk835k/lVQGkbkxbL5MPQhoyeeJEE3BebsdkNy7UZJuhRbm4xljIvMNv4h
wKv7eKHcNFXphkqEA1mCujbg5VzMsEXEyFO1zyvZ0MF51GCF5qrACT4qSGjY9KPavO7jLsUTKxbY
B7nburtBmnHlZ27LP8jlt2gZfJRjp5vA+ihB62OFvATquWvIuQEP7tDp08pQ/Nb0cVGphUXYiMHj
TJauI/8VxzkkA+ZdF5GaiJLbBirdG4wg+HR8CkwgIbzvHG2hKgJQRKJMDKLgWaDSQpDjGAbn9a/a
evw3nXAKl30DSWcZALnxAzGbrNFrhYhkHzahJzfifxQWr6u0Uf8aap8n+DF/Yn+IbCx6k2a5J9TL
ukZ1c402hbYwTvrRg3R2eax3nuG4hD1Yzbrj5mnaXIx/IQZCkRFc3kkJx4mlsV+O4Uo5FH2VMP2W
oX7IYt3pJWSbGrMhC4ok0Ic6ikx8m6QfRXanIjZ5fy+u6YYu+Te0LpROfrVM4FCZZa5PHIhk1w+l
S1P1hplYyNpfhilwo+wa1DaTWnjfVhl8vr/hDUtraOAurSkYg2mBE5WmtdQeKiGG4x6UqwEkIRPM
LO0JGEhnvVHhgZtyIiAwMJcJPJLJdV/7Qz5QnvPWQ7WFdRWFjtPzv5MFnJkcSvJMzCwgGGl9cPTD
jCH1qifINsOMHxtK4B0bEbHlZ77RbRrCFZftFhdL8E8jN8jbv2Cn8PL42GVKRi3NKZg1g4/TJrNe
8+xKNXZxm1+y2iv1RSdlL+s5oYrKa7nQH0oOQl9OWRRgDuPWWw8QXBR2wtVYZKeLUjsu+qP58HWQ
kO67oxG14bxHAqVTjmg1lbmrJBHN9yRICx+WEa9XZDhGMLvpGE+kMxbqE6DhSV2/QeHqFWea0xk+
X8ItLrDf0N4QXbKoWM2U12sfSLOrhcErPbk0wubNc+pIvVnebGHuh3xknnFgrWnmoOrC8nDIDcTk
4paoMueXZ+5JtziqlBRVUjgyRZI5i0KCleIEjk3c8Jkd6vo/7HvVgqAICup+dlr+fnXtlxHkzbZ7
aBDA3x1tNBfiHr03N2gd3bvEWtZ41MKE4Z1NQtl1hHk9ZMcHy31+ikQnk1lnF8Bt7GXEnTBP6IbB
IjD7jzbzoX22h7zCqttoVKBp4uNEhM+JX7tS+QpGTy83/ScihOe26B+zCa14G2/yE0+22jP2YkOZ
sd0rdQbSXs5EqiCdyvo/5YxbVQLkLPYL/vplvozeWc6T417Gt0agTI/r4wLk/m4jYAR9TbBsc/Pb
F07/HcxCorQl496nNMjl/q01hs3qn9RA4MhJFYpApAUTT/VQS4gLUcG1IGujRSjkIuZ5LGi3UlSw
qUhZEdbX4rFEfFvb5P2VbbNvCSgJ4dUeNLfcGwAXhhIe0KnabBexWmeZAzcYU7ncZH0DfjfX/qmn
dfhA/W8tyXv+jUHIkuzFnTArCF4qVBT5ijSpjOMBGDy6eJvkhhma3jpSOR7JHXi3TGziqZCn577I
ZbfpoBtJaiytBtrFLKy4ST5iRo5AJFMcfyXcS9s+zRw3vV1yqVPk2ki6LJfxM6TlH/bkNTm8OsRR
MqPKQq7R2QMC0IHs1bamTh9jWbBwnVixyceiktCD4q9XX3IJlJyGOr7kowz+cHsTDh3sU9XoWJPh
5O/sIocUN6dvVftgme+DqlC53T8CiimSsQENsP35iah+jeYK/1fjM3Kf+TVi3yRwT0d0HMJFAg79
3vsjgYSSIn1XFKOhNMYyhThxXVBUJbutKK+mdpwtrIly9To10H62gLdubYPPHXfR7ClE2YWBnVsJ
rb5DW3gzFTgF449V4X46o6MMZJ+M2hhVXlTRsZH59eoLXzaBHcJZ+/DowT3jcYnSKvWi7fQeqDC6
klTqcp4rx4/n7mS3OUKy+rIKr2SiQnAtqtldvaBovFBzk4x59dx/DAFxOeDXcP5wL5Dt9B6dIj8U
/e4GVWXr2HEA88tbab4KF0NUptuwQ+XYbqDziVqTYrpatVnJecmvo91HaAleRUnnM3qcohfOaeIW
t3/g6ByBINXJN83Ft1DdYXGkKHbN2GJDBgu+Uv14xz/seszCUQtLWFq3tJJaWhGe/FqRsZOw/Kpj
IZd3iruQnfUro9ngMFIgcts8CC2vWwzlV9Zzi/VJd5RZtJEyHtP4kd2lllDwyAg+aWNUDgZGQlUc
PsyhQQZ6r0Y2r07ezM692tLrQxlBpqR86pALUQWFgkpW1BgCC63zUnvIzpK95h1g/gcltq77mGxx
2esEOgLzgwSNfhn8JcUnnoGOMfnGDDk6SoOidSNcY3A7ZJ9fmAusDGMVoIzg/5zhY53vLsYkcUlT
buAtFNSqt89S3wamyD+Q1WK/erwNA/pwfG5gETJnd8hxMU9AGPCJNfKp5Rd5mA1dEImqoiCHceJX
0dp6QHMaA89aJxKvnmkM/tzTR2PkXeEEDW24tWsiJjHCzVX666GGn/X0kyx27B5hQwICVJvKSZn7
64d+yTeA21L/++tYDVlbwDrJAq+lfYPEMcFJf1l6Se1x30Z0za0o0bywrfnKejKc4KEcFetObOVL
6I/au3d/Mg2ofwEgQJQhjSUsQdZHi7sk5XvrlSbcKwX1OcnO4bWfBybBTrCIbGUz56MBWrPmqRdO
Ldah4DHRulCDKiH+jtfQWmMU9ed/pPY5Adw/CM3zc2lsCLjqArqFIWRfEsw3vJhN64nUdl0bEqtL
+bZqqhJIL/OghqLQg92ObypTgtkzUA7pUXWG0T77RAmnAAncEtrRzG3t7mV4qdCoWC7Qj2miSUJt
M72N+7YPj2BI5i7HoIDNlpPmZGmQZUhy/Lsvy9rC0OqHn6Moh7RYfjKFFS2eHuhxqIx1G3iEm1Br
Q4VG3qPPvORTeDztGxsuR1gZJBflBIIo04C1+pK4QWDm65Mn3ZSJI7Dthue/1b2XIkAmNQPi8Wmp
Mfzz3aH7XosHnhGzF4KH8oGcWjXk9GSE1B4hpORz29uoiNd1BCAKZqbF3kiho1dp7RsZNl2bk51m
n81nC85ivBSmZzVOjDGzlZyORBzaR0OTRB3/lVbgLek8dUUdjZz8HsF5AYfhUlL0F6rvC5hXfkeE
qw0GHMIxD8mcNjbnvRSil/prJQ0N8qpazhH5SYtkF6ZZLs+yf2HHFZFRRtO3uZ8ChRtaeooLByTO
SJXjwUB5CYOZo9lBv1c2I5hxfUqOVJobn41z3mtNVcKGi+6Vb1FPJ2AUr8W+Eq3z+xYbILOdasV+
a+fBcXXloCSZej8hil6fviMpxhQ8Zr/FSkfUJWFyYoxIiB7hQ9Q7bstyafYENtWWJXeq+9yvqpgQ
nKz3cUpawWEAT55oq+nUh0Ju+oBQKtyObDjIYCvpUEJD3pnMgnCFDiMOyzCo/CTQknMJ7fG82ery
qFj5xlTkUHQaW5BqqMn2aPIyTne+vL0QOEeEMq0QrV6QlU8uyViLakr1YWNAvQSisxJN/NzYEkI/
Vwwotmq/KoJrIdadwiDiIixCoIZFyDwHcJ3lL1SkIrHLwJKjG76UpBwVmqYlzBYCpwV6SDUCbvoD
/jXbSyhRWXmxdlLL565uOymTMb13pT3jU1vRv76PXvPdiOBUWTB94Xu4/A5RoHL7xEoS+Ida6vtg
rw2NbB6gXeFd27Qtw7npkkjfjKADWNFMfq+d49cbWWAMPlEllkKapixgqLnFjIGEFr7ZwK40j3KM
zVaxCly4nj0NV5AMPsbhrLfOgHpPe22bi/xz9SsXkwP0WOIp6Qp3WQfaINOtjq6xpDrAxuDB9Ppc
Ul+W/WIg3/WGMHUDx354FNjWVOgBE3uRdCLbMZkVbbZIEBwJ4sPX05kSg0FlyT4lU71ujMe1dFNP
6R29iIeTuI3Q0sIz1pFHu1t/IrWs13jPOaI9uhK1hRrwUzclp9jVkdubRocaLyyTRGJy2UHLFpQ9
QBFnDGRdwhIPY7jK3IzyGfVWJKcpxyqg1CmAfwRyEAnOQWRC8KBbPAv4OE8bAJe9Ew0h0rqQ1lfh
lEEaVwnRpvsoIZDh2850ppVpz1zs7OreG1fRMiFSJmtT31gDnJ0EC7EMYMmWXrXRwaZrCIui6UCB
zmdXhqQhrn1r5Lz1LBJkSBq5nSu3Co4QgUi8dVwkIhORXZcx5JxRh7x/Su6++w7+4g44evFjEwKO
2fzrExp8emfrXAeU6uYjvai+1A/GiF5YX7qeW6PbvtUTkzCllOuwihOWRrm1JM75pNfi8uskEHg4
CtW98kHy/iQiO88PrqKFHZQlDM30gnI2mec48Ti7EztDep5dxApkX+9OIwwp8BiaY9V7Tyhup/kD
HXL8XANn/GTDTpWGR1bS2qvRvQBFaMLLuEusWskK4k2NuV+q+AxOpdCn/vQSmHHFjOGf5/1zG6rl
rufJFpSX9rz9aE2PItP48fH3T8Kxlx3gPBPTnVNv+2jnsrMiwBXeVrFGUy3hjDvBjH5tZahcUH3x
AIzNxSr/m8Bgbv0SsQkAU7olWEY2Jt4aJHJV1CnZP5p05iRwRPmMppNcJi5zIlGL9QlEr4YOzLeY
w6EZCMeod61E5xdZ9HR5ODOoDgQlbqYneGjhp3fimFwI0ijzJrIOF9zwfXoJDjHf2qyTakvHL2wY
s0EDgxtXFd+nNVFVX6M2sDTTXiLh/s+yh/+tsuxtiayZWkvCL/BTO3o1HCbZd6eV77GX+3T5PO5i
m5cDg5uZTLYKlFPvK07tRzfnxVPZ7ZMzW0AnL4h5YlYeEHRNHhhJ+mRwIU9Xjx1wIujeB0UA427W
wsOkxaJQRcA4pMvCAzDoxLrlUVPIrz76xbscup8YBYPp8NC7277pM918cDQPchV/o2no3fCezpKf
7HCzB8VzSWeRwljE53GrjzNLBOow90GhYHmLAu+29Fy2H5mLG8ERsdHUAchgOejDtFC8pVRvx3xf
dN+pd5P1iyugXR2YGT5tgAruGl0mq+LzbBM1L1HGytEQi8PD8SXZYe/SZiyxM5rbemRaipHpD7uL
sRTLUHBWXt/XjPeqy6okic9MeeoQrbq9kaiLYlFIVbOApeJm+K57G0si4nz3/nYZvbOTml+V+ApL
uO/H1nWeKHPBPu3XtBJNu4QXmXkJuRmJ//PFR6PC0ZIQES/0u/tPPyGz4JdQAYECXQ1fuMN9Q7pm
rdr1PdUJpJPzWgZNDmuOP0VqF158Gy7GRFu3iPZq+izwV93268d7QtXbVE5C7IuLG4IouHXh4Rok
pZLQjVAby+RHSv03lE5xo4KnLmS0q1fmQKvyJnjRuLWzn4LcvgCEZpvTFVWM6LZo7KMlqZwZm7YR
3jEvPwg1fjsexr0Iev08RI9qM9H9o9xLhTPkRIL/ziveHzSOVC2HKAO0ji+uVDcRo4Em3nswftc+
fWUj/znZDphIVa70oh9nKsY0bl4a743WskCEMV8yaYYo2F8iKnXRqkRdHWrBvvlHQM6zVWo5QjGu
UQOlUCzKlb1vo1Om/nStoMXLcOGwI6c35fRxQFr6s3lZfiDEUic42yV0TWcLFyZj8DMgxgNJzAzP
EoLgbnpE3HfojElwhKoCSCVtxz5e7ukSpzU5ZvcX3m9bUUjNthi1YjziI6n2BGxSE+Mh3ciskpGC
Zer3H/rsI4AB50EwcMyOCXQSIA8tEN3Kc+3Acne60zHcEg1XGLj7E5naWxq7tWxz8Kvm9ZQoS4/1
a2YoZAKHwx0nTByXfVz1nEXpSiZP06QJsMmXorgddjpDUHSDcSz1KjgrsiGNL+718MpHqiCTEUIs
10g1Tcp5eo9brLZYGisblCKneGYsb1S5AXNysL+6iqZFLq82GqUGQb3GgtLzMPhM7jKZkQEYs8aU
bhiAJLwaj6jVzBY3zGsDWZfRmN+bVnqOYv0iDdVypgUFR7AgkoGqC/6F0wSKHf0QZGwYC+rXvOUv
Ds7cFUBOcdb6PQlQjZGrADXL4FlupN4SaZ4t1YHLrfd4EHq15w+mGSNj48mwKeT+KWT0UhR1ruKk
pJQkUb64It9+2VPnrGLQbxp5m1CBR/+yjYV3OfUaJWkRdpcJlYnU1+irtwcWsvIxGTZIrqnQWOja
gqFqYVn/e7fRDbleJ3B3nCgTMLw9rL58H9A58cwal87ctXANNCS0HM1qouf6RKP0naXQjsNc0GNF
O1b+E+LL3JwTm/sKj/awv5bEYGfzIVlNfpggFcO3OLP2smwy/C2P916aCMU4DDrddNB7aUZwc5dY
FF2gAH3Z1K3qJp7DbCDByazfrDC+S9R4GieO42FjDnw23Z5aJ+9Pqc8njvsmTlYbdU2PJO/H9VNB
IVoM92jkwaoynLmvefdbHDyqnINamV2jqSqnrSWjPMe9ALHwpiH0VfSII77MOsUeUoMuvEMAyfl2
4hTFLf2Xqiy256jNd1a5mwIiPyBLDJWNloyhBtTDWHojnDkw2dKSQZqSIaiFH4yIU2EI+mTnYN7L
UH6tbWN2yxFr+L0PKulpYB7IgebaVcPs5MXTekehJNIyD5Kzgx+ZyKUu4xRx03MjiLN2rPLU5onj
cDBrUhWKZjSx/jZW7iQWI08ZD4DOMwkFZe7L1SnrYw7C7nf2NGJHri9vpwaXmZRrzVCPlno36iTT
/YoVJbBfbF4JafumJDRTSErP4Xdl10EF5oulQ0RVi0MJQ6+HXwHLfQV/KvMbc0jgWK6F8a5msDZw
TJpZR/WNgsVS/g8ZAgBw/ygAYhFBHpaDckUH9U08N6h+6kHq5trQ9WvxhkbldOALkWumG9XIDWku
bvGouriB9Yj3xbiK22sSSK6AnMdfN9m/WXorFsaziHaH2csJ+aBAXgfOh1tM4zhiUgaCHHxzRW7u
p0DMwoknqSg4oL7M615x5LC0R77lG+bPoTlrEPXgoAsTfLcv6MX2oPWmJLtxVgxSaQjb9Dp8+Jca
T0uVFNo8eLj07DWw3Ewprb/8RIBnDXe1v1Mwptl27EOH8pBCaSeNV9J8Jzc04e2EfEd3MB4RuCj1
ROSMc/YnDLubByJGXy/rUROUBLsDp6usKCSGJ9BmRoltas/AzOTv3WaoaJBvUptWE8midT6mB06m
W+KscwfYT2LXDx8DhLcY90yr/HmWETGF8bNRqy9HlqnneXaqktOt8U+VJbZUlzL1RohDajXkFkXA
wf6zluz6/duNsfkJM0PwvDmFJGTwOOkFQLaNcSYGyNq0prB5drPOHfkBXJeM8mK1f2ALxV1g9eGB
tRaDsb7b3GAwk2E3kYc06wp+hU/RkRESwXA+jpyVa7UlDpd3JNhY1GxER3TxiizyCRXC9oIjm0Yw
1DwhgOnV9nPeX2WW//qPYJ1OprI12LXGMZNkVw8y1YtgsbfqGO5HiBjG2E3/KNF6q45IQcav94iP
R8aeaMdCxZR0rXBaGlZxwAYb167stkunvu1qVjwxIZiHknoM/2gKyTIZR2WVKM7b/38OtbclPXee
Y/r5bM1WOpaXPwJuGN+JtMdDpfj/KkEiGrpSMNLFoHvFmR1AVa75Nq5Agl8md7bMuBInf+0/XO4X
9h2Y/0236jpaBlb9n0ID3fZmYqojIFcVtOaru1KnD7MwgumtRlso6mF2JsesP4yCS4D1Bb8T4O4b
45EzM/btWddyL9aIboBpqGU3GAqvg7fmOSpMnyGJM5KDVnrKnEv9jpBNIVZbiQAOrALp+X2Y3Bg1
ew7oW5RT9DPCExQsnW5TA1AE5E/TKrzP6fjo5QZVQKoasD2c+pR1YYYrP9JEj6o7VPabKi4aAscV
wtj2xQzyZrMuDO8Yr4SstpkGQJ0uCaRKFg1jlo2m6aKIdz5ydxzSofym1O/tcgjfd4PG2XOlBkGw
q7WwSvl0rvKeun/0MIx7IL+ZlceUOfbpc4Msq5OoLyPU1lw9InZpd7ybo0nCaG//8h+2ilyqBIVa
7CqA0bIPZFxbIdhz14fxuhBwUvAmnk4VGrnDR0IE/OAAl5BE79IqUKnvigLPfLF/vK9SkBH5eG4d
w16drXInUKYqmI6ej9iHDfS/0cgTDH7CjvgaMjOqh+TFcQRR5MxEOsxR8g3/0+C4173BUVtSYLUA
Zsd1eXlhgwclxuB9xY70UxwEQ+5D8HrnHipqvDpB/EsWat0sxXNjIHfxUWlDgMlQdSWjSsqN4EtS
U46taesXp/3/aFVqznTCj+ZRSqc+9UZ0KO1UTmzDHR15BTgNhRP2kpQjeltkwNy2thKns/xLEbMy
Vj0YXhNJdMl9xMnWfFV8uSjoE0KKQKbepJBczDiGqkyFx54t4uskTeXHyJba97AFhbn61b0bz+hq
Otl7Ni1rcB/FTX/bag+wmTa4Wy2KgN/4GY+A629dCCitsxSbz5lHRY9sr5R1KvtZweWcKclgsaW6
1HVzx0zGXm76EP6Qlsk6hgJUiO3yxzo+ob/BWhPmbYeOG8f9AxIwLG7lmmwnHW9LLvd/hm48Obqm
MzSKR8Di7n4KPm5FNBsqbHdxX1VwVOQu7g0koX3TuIqsMgBrLJIztFyQTC7qEUR6LErhKOT+Q/7U
T5kU2nhlNA6fMhKfPbR9sEwMkkzMy35L7d3P5iyyZgbmT06uJVU53nHFhKuxQyafgApy9M9MC6+f
eJ4kJYaxrMUbnVSIa4uH/ba1VVNOWg2/XzGHuK0SVi1wQlbnQqy2dbwnqaZNeJH6XVM+z9kJ4XSp
u/ubCwKG340yaWnHjG0TqriA9niRUfBRDATdTQI2HbqzEGMd86YqAEVDCB5Jo7XEoBWTLZglnnAi
j0lEX32P9QL4CLtcfKn3pRykGWxZqJuog/ljE/6r6wswQBRY/9DwQSuAtGGDDTuI4vm5G1977mQZ
eIBZ8pezJ7+jH+mZnQcXgz8lQwNoh3K+I5/2ziKtALzE4xlenZidp2r2/UvsBVuSt0dkNfZqcDVp
qPjDj2vKTmk7w1v7xlsf63BG43QmJYp7aoZnUbT/WL1nTYYlBEKWnbt3E7NlIDnuZTTM97iECy6N
8FZlN6pHPKtqe8ct9HiZqUqu1SjYgLMb1h0ggBDHDQoDZ7nm55Fkk4DJdjJvS3tN/TecchcF5+pA
ufmYI3GX/DikiJtt15aFn7p6GmNKZ1jiB++3YEyJVrPIyZXsUC7TVIyWeVQytuT1UrK7i2s/Zjjq
VDRjicUTVR3lLkDU9hqduIBIL68N4i1XrB5IB/XyOZL77jlouYhGsX76ffeLwVX8wYBZLZwvm+q6
YX9ouA6oNCWOQi0mybKR3o7x+dEFuw9ysPtYjTMUBHmHM7S2A4Sf7GQr3H+a60Y7vfdTu/+TLGfW
JT1JUS0Dw+haIBHgwXX2Drf+SIiLlGNXR/mcMiFszYM1eKYNnreSjTtGgbrmazuZVROckIitPuJ0
hKV54hCH2i8962bmRSr+Hyf1uIh1/h99HSTw3w7G0gKfQkkvFD3F7F4DyChJ5azb4rGyuqi7biuU
MzrPKf18o8c/znH0P2yILB6WN+MZ5CMGC4rHwBe+nY+K2aNzt+/UD5PJcCy2TvoR8fU3K+e6e4r6
6BGxxc97jknQml2c8lwATf0HWMxVYaltK0sXFMpT6jcTYJiZqdw+DD+vbT7bgAaUMcAjPaNi+shL
VVXGU337ZzVBI4neVhxUtePIc2uYC6RI2C2qxQgjPQ/GTxswx7ukdclhAv5bVRZCD+oI01UD1bEK
1H0HSpsdor/2iZkWE0stpI0A5C48GubGM0ey+fVXcon/R5VwhWcj5ZKqD3S4TotmMZsZTdS5BAv6
rK9foBXUWUWTW5rJ5Jbhb+WFOuIzR+lBUOmYAb3viV5P8O6lMchOjqWpAr+v91c6KOksm9hzBQvw
CcGi4a6tdwGWjrtevguSbLbA2SROsAt5o/8VI5MS4kIk3cJ4Py9UWprXtloPLHjuX1zPZkOYlm2E
6XUzGYjS7fbIVXOXGyR6Y4jAryE9vLB0Qv/LkvPLwLqFPG8NDRIipNOPuksJruUhweLri2QmShS/
9K/hWhrBPNyNkVu9N0yjCS0QfOsckZOzngczFcv6V/r7Uf/Jobm4NbaKs5FO/u2BBToJfbANLSGV
+DG/BN+2iI7tYoAf9vdIG82UIWM97fWDq8Eom36KgPbQTc63gYfjU0KuRkZF1yLRl9bemqAFeT7L
rx3IFsKKtkz0P96lm0yS1cWJQHSUKO3tddxUgG87iOpOAFYAjOefZleEOjZp8Up0RlSjoN6CLEuz
/Aqdv33jOgD4AUivP8dFlNwGCjTOszyeioMZ4YHZtOpzGS9RFw3uqo8rKwfR4S/7bAElAUcBBQD8
MT8hfn/UifJtCZ/udePcmT6HW1oEwxI67bwQA9gUm/hboXEQoTep62VAz5/v/boTpwGS2KZep3eA
adSeO2AyMi7WUgjSV7AE2G/J8+quZSVrlYM0H1yOa656enOOH9Wy03pMqfGEoUI4oO5lv121YEa+
TEInuon6KLBGuVhqeFvky8JPfF1GeSdizml/4iSvY5/uV+RMyLLaohzptEWomu63MYa2GQzCtbrm
5+p33cJVkSNNIWOaH7dGpuvKRhBTegNpwbBu0vRexQK5JFFn/fRf9cj87oHYzjgkIv6jvN2fn9a7
W5u361M9ijVmoBEHabJc5DryC5bdM2FL8KtKRYz8zbyIzoDoHOmfRabnCw26J5Qczl+KpWMk4nsd
1ClBIcgxTfcxnN25k39bBVgRcbkNLnwCSSS/4/DxOdLenCtPVB0mvMVQ0+egARkSiDKvSan2e8wk
ipMwSUUwf9TDzllq/MX7Z+bu5smsvY7Q+fm9s4cF4jXqboShjCVu/6YmGi9NBuQ7gSdMwRgCQ8Z+
GuKUm/SsL8wdCgX8+31srVzV1FivFGCoR2w4jnxy74wWFb3qB6M80SzSrN7C8C8lV1sr8B/MZ2ov
EIjpKiu9QWm5ZjyZ1jRVJQFDbQ1pOPLVGMYz7E7ZLgX2bCzBV9wekY4299uOq+A1mgJwaP6wRFsy
C5PJNvQ6E1YoIGifyQVEuC6ygAA4UHkL6iJTPQbNXIA1QGjyMnJODZbccvagm3OftYCnQqbyCY+D
XTQwLsA4ChnAI5R0V4tkKAJhpTF8zmKrNxuWzp+9fwimx/iiZGjZ/3ghObI74RpnZFmtwA4a0Va7
2ffNj8MxSyA+vDn60IQ746CVQm0MisfNkxOHhm3eYqn4uX6QbPC3G1z/8gg/8eDbdtzLJKfDeRBm
mCGJWlkOKa2CIxiJ75bHj+f5N1v43uAkTPSOsCv3rnjGrs+TNQ124mmsLppy9QLzIC3wRjC8EMbB
NlanOREd6ThCrmlADlAbdRCn3/YaNhw+fdwGfnf7Nd+69O5NfNqVsU6ntRL6Icg9vC0HsQSPcFYy
/asCXs/PnCLJvVfpyMgRRcF3cu0NeqsQ+SsUjvmuiU2UeygNlkhA4lOKOmRKQa8l/LG0qJ25RaQl
KfopfKyKA8F7ENGBwewAreAZI5LT8KQj51YM2OWXOmXkhTf2IfLNX9Ost0Y02s7YbG3UYQCN+CQ0
jT1VpxIXOlpPfMSDY0G7y3E5ktrblITuJf19Bh23xsa5M9JUYFS2OGS443B+ujKirl5Vu/+gW9HR
Oos1JgqIMbwBeSqidHdXlHYzJJUJ6JI24lh0dzUztYB8sCL5HlMT4GXbDnamOULaqpyVC5nJjuXW
h70gpVkR5BvXKbzSEWBwPDNF1S67JyJ4sWZkcyZ/0hGiwp4kspRrMyY2vpKCYPOwB2P/rXkDA8PP
l9QPCB4TjXnnJIGjYAsEa/k0mc8XLyxk822seugpcmpdI3HMjwHlO2gHtUVVhLeVkTB7k0+0kdae
HzSYUuVM0nt5jIlW0CtsNtIq38dKQ6kdWFhwXbTQntslfh9rohTR8cZMJo0uqnKs/2t9I7qYIO6v
ZD67LyeXWo9G6iA55nDMl4zmwF1voHBeTEEH1nS7tJq2PEcd+PwBlUk+4iTUrfwZkay9/Gq31mOT
Ybctvy6GI6l5jO7Eh4sPxpkRS0Wy1uCdTyh+SURmHJpTYzcnWqxwt3+EYi1R2oIDIJO91sZhTl08
u/hdIIb/BEi+LJvq9REcLEID4aBqVQ3slAZTFP8MrkcgxYUGZ+mU44LYzZL56YNAk5gTpGuulycs
ySFzbqRJvHjbuX4dc+20G/F92JYqaG4EzoSQumT8p1ay6BoE5BPQyFoy3lv4vrpNAGN6kRLKNHyI
6Rw3ZKQmxSyNcol4iJauSab1FBvRf3LiRmZAN7cwmKFJI1Rdlr6bzePDYW48u1vo+HFQNh2r9nyj
J48EYN161lzbUZFdbOqPBwRNKf91ltf4mFIyR8CwN3TkvsSACPZ7RMT4/N4ywzZs/SPf7O1t2Zso
tjMI9VUW++fNArLuD/MDLLr0aPXUc+GTtjX5wFrMtBs2kIdGgVDC2N4LhyZ9TaM4AKJXFuI6NKcZ
2lScSqT9rfz6Af8jlrpcNnB9i21TOZ+HdAFC5Ys3cCd+QgSvIlBZwjhjdkPx5aw3BvW7+0+86IDE
VEu846UycPpdMmt34SyxBHpkrfs3EUQHnJtYM22HvD9Mno24V668B7o4L3RCKMgp5CN38B9hW5tU
54fsT6tU6LokoTY0/ueiAbmld7+kgyrsqtLT7xsvsLIHWu8xnqoJmB/YT4lDYMruCbkuLQtLLNw7
yWjO1SL9aMgSoT/MUioCMHS1/6SEXLtEKKUluhlCwv0DW2pDbirxwvfzjkmKvGmgV7mNvzMxL9KC
7tHeP/ZxMPRwMm4ywC6v6JcYRLjw3hh2HZXDBFmBK3N5NVX021vp3oCT+YvyjbyNlK9Xr7GG9jju
Kx3y+2+KYy23kLY3hu7xEckuT0IRz3upOXrQMd7IJZu9xkOJYdiG8MNVhxPjvS8a9GExD+k0h/RK
5OhEVox92NAFXn8YGSwrYKfyMH4KxiXUqlIR6MIBy2/NZozC8rxR8sCnCDl9lezHruE3JSV4ZmRi
9pk8oNu6oMVdRcepwi2CRLLnO6ZbkYwlG6z5mAHq/bzNDEjkHm8Zf6DzmNR8KameV9XAXGp0MsyQ
ev0Sj8UZys9ICJu7l2ycNq5ndEalGfAI3ZMII2ep9MgeJJMcfqSEvXzqvRnOFq/vKTWHTNKd3Lby
ko/MgNcdwe6jwZMMwAi7cwjInbbNO0/bvfm1aguLzvDVHj7+zWG7QpyI7Sb8diotAY1zk09TvrEf
MNLte4/ThP14r+zCSq4x13l/qFSe1EcoChxlzAzlFlc5U5Vs5AdsWzw0XUAnuCdC75DFfsiepWVH
rV8I/4Fi9FJ8iughiAbpCby1kGiGCqxtlu+WhVF3pBi1WvCTjUMcARCP3EJKMW1BQ0WewgeuHeEb
x5K8CiHCtooBU2+yulY/JraRxo+QPZpSS5lA7IbCYRx1rDlGmQN5pf3R2sTmf61SOxGb5D7rFpHn
hjFknMzOauDvEY73UYRyOz2I+O99vDWtA0yU1XA5lIz8E5zNuLEVb7S1r1RF1A2iYwIYkX4JmLhE
HwDFLbOvD8FHYgtLo+UE0/qa/6QBussyIGcWfxwL1TmP84axO60bPueNbNA9dH59ankiRu6pN6MX
lpR/Er1EI5iziJE/8Cqb9ofukTTOHle+GxQHxlNPKoCs/Or0cW8PPp3E6Wst4W7c0RjK6FDGI1tY
QOVai997cfmK9E8QNnKnBbMDuYncM8I89ktGcskkeqD8zwYHudrDeG+vFIhGbTwTCfEapzoCSw3Y
4VQkMehELTjBZgGMTtc1pXVLKXxmC+ZRK3iREjQkdpbaRKT2JNpUVVTusPfVuh0viFm5/nh/mk3E
bwWgQAhdci4XuEsweduTmBz4uPkRLCRcBbqPm06lsHX8RIkTzLL4F8pAlubQeZxOsLwak4TF6oqA
v0Co8SG//oJ3mkC+7zqhuhaFsVE5OWcVLmnO+KpJIqF5FEZLlVzsplrMyr/pEOrGR4MKOJRZIdg7
lMi6Q+3RFMLnKlmh0X2yNctClSssN5npNR+7L9EJurCkm1WAnIszQQx7oF7sFi3Yyqd1Smwp1RWB
WkjiZm1aCQtLdrLUzgtKmyAPyDLun1W3HlA5AWLAGDvI7NW14vI348v4bRDMNh737WcdUeNCqBKo
5Z4RQEZ2zNTSA43fTxzaZT+ulbCVEegl+D/TJ9V3vpeFlkuR4Gh2iHe29gXKbcfd6CPuooAE4EfH
DS40iDMtc5b7qBrgEVUw3G9nVzaEcvX2Wdd9f+ukXHQEEL2tudqVmOo2mmITj3Muha4yWnh46KRS
airuTf4shze9BICycepZ7YLUovWU9+JBxSynHQRH8l7vjnWIHDcIjjj5d+bFBcjK0umZcD2KrESe
uea2Zb9J/1HYZbjMSlzuVK2h5OLII4aYWmkjCCRqiz6avGgHWmxIykM8G58Cn8WQaOijlgs5/mb5
YEEzB9ZeVVzyBlUgTBf3td4QBLNqaYqDEyY7kfa2erg8UyAKp6haVErmQ26XrllpfXOPKQPtmSvk
Z9tOQJ4DLX9n+bAKnmw2+7eB3TsnhR2HEhPKForC2qkSE1GDpoSOjB8=
`protect end_protected
