��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����N~@#�k�0!����+��=L���0�ԴZ�2�Mc���ZO�����=�����վ�	"cqw��a��TS[��{=:�����K��-�մ�(��k��N�-� 偙O��QZ��~rL'�x[�i,mׇp���O�I43��4d�,�H�����SN��d���3���r��m���̨T�I;uj2Y� Er�*p�Q$Gm���p�V�`�2^���,hz�<p��l�Bxt�5��s��\yq���#�@W���f:m��T�	,*�񞭋����_��㧋l�	�\�:��uGd��PǷ��N�I��_����Tuv� ���us�(H�~�{2H�:Zor�Q	#%�3ˠ!��iS��95�,?�.���/�F�i{#���Tp5����Ҥ0{%���2vpn���X�����@l����3dc�ק�3	�Ed&3�ZN O���z��s�yxӡt��v*}ԫy nj#��lc��m戭k[��5)�A#�����8�!�]�Z�s�M���t��w�!��'ÒE�rv��Ϝ�c@<U��\tq+��&|�&X1)C�����r�A~��B�&�����s�:n{p��͠R�X⺂L^��R����c���f��J^?��ܣR�O 1�rV���:��T�4���AD����˩�F�w��)Dm�O�b,�a���1$��c��7t[i2>�ޔ0,S���󧇳Ϟ�ᒨ�-��}�!6��Jyv�醊�^_�(�H�(y^����o#����X��3-�k\8�M�T�"`R�DF6ȕ� �,5�;Ҭ C�k���1\������k�t־9�}���� ���QHF��"��t�9 ?��{E_�7��!����](�S��0�q��w�9��=�i]�1�GʦȪc�W�XC�|�$��}q�6����zf(����լml�dz������*�eLD�*�,�m�]ہ6����D�Gw� �g��' A��)�m���b�����L~�B�3A�/15�s�dm�\��rbY�6�g��x��E����Uf��)
^fd���YaŌF�<����^ڍ�-�L�A�hm�Z���JA�&�拏Ӻ�*�=�#��Po��[U�Ƞ���>�-:NM�)��Μ&�^[\c�s�.��i�����+�G'Y�h�8�|��d�j�?v�,�e�Qy6p#��w%�J������q�O�U�>�(zHO�r%�`V<�Q�O�+�Y"��9���1����zlP�
�#�i7`Vq
|F�L�-��x w�lP�)KG�m1�V�Zq�����"�����?1r�hm�?L,?ɻ����c���6ғ��#$��a4S#�G,U,��^� _�&��K�n�q�%Р6x��h��PXL$�	s$m0jJ5��D���G�V�ss��6,H�R6DWA�����^b�ZСi�X�����0�#Z�o#W!ZH�CW4Q� [��]Uq�%}��_�f���������%kY&~*��|d���)�O�/~�#2k��!�����(�8O!�K���d��̿���ї_�5Ӌi-amC>�,�PF�H���uu�!�`$�4_���6֤�}��.Oa�f���H�H����x��O�Nbs��r�|��k
��%��g |tHե��b�`#(�s�ؤ�[X^��|�we߃�^�~���)�y�9Ӣ(n: ���������a6Ki�9p�Y`d��Pnc�F߄(����	�=��޿��K8.���_(�b2�J'd�o��T� 禩���8�;�)��h���S+d�IyԳ�M��%8߆�8�?��$��u��:�~�f_p��K�_�2���7K�}}����h��|�U�5�@*�Q�1�'OٰI�^ƴ[�<O����>:�zF��!¡Y}Ed�yN�.@���D*0���?]�م�a���E��9��wD���@�Ԭ����g�<ɦ�i��7�g~IN?��fR�WM��5~Fq��؋5�P�zC�6`����u�-g.x3�,�sYļD���0���M_,|��08�7��G�VY�f)��n�MZ�6dAu�|1�&k��آ(�%+�{��$���כ�@��_s��Q������H�w�����;�VCE4o���� {��׏�V�i�9�U�S{ɺ�
����4���	���s�	���c^KlQ��>Vz���]ƙ�yTD	k�����5c���M�6rw������U@7�-�Ⱑ/>8_�,�GF�����_��ܳ��t�����U�,.a?<4tMG9Ҁ�N?��;�Y�v�&��}�Di�'�u��f�U��\�z�t�*��\�f̝����B8���[����@�;Y��j[mu[2�q�'���F��r�'^H�
�(!�$d�#�ʩ�-�{�5�E����:��';�̈�۷�m,��&�E#�����A�ہ��5F`vҲ��߭_�sm��L�k襣H>�(ZsȈAF.a͋����jD�TEyD"����U�5���
�r��L�p5�3�����-�&/���x+g�ވ��v��Qzv.Ѷޒހ
��s��V���g�VUW���;g�0R�צ]3A��p�D\T��=�6b�q�u��# ����F��]� ��KdI����ыC����籆L���7�S�,W��֣HF<�\�ͭT_"� �"��*^��&��|�=���*9�T�kKЯe��Im(�ʞq��t�^�_-u�μ�\����>	\��e?� '遟u���G���kn�@�T��i@�|����Ꟶ�"���U��t��톀�X�X���j'Sh�{�*y|{��}0S4���;� �쑵Rslә8�-��[��@�PDw��]���M��G$��?T٘U�h�@-s`H>7��ZЍK��T˪�a@L�Dx
uSײ-�-}̈m��M�r���;��c�Wx��M=��O��9��	a�N�=<HG��:K���������+%�N��K�]|>�������nMXFh:"�v�5��3���V�����b��R���}˫�2g�F��|:�i���*�jt�A�-�U&������8K�W�opS�tN'!i_�XQ�ڀ�����@zé��0��椐�^��j�Prr͌�J\+��a+�A�X�3����-8�:eR�~L;v2�Z)~�e+���֙ �v�f�zoO�n���0;b��(�(=��Ug>-gZz~�>I������x~���U>v����GeA�L}4���8l�zz����5�3θ3����S)	� Q���sS��{�?,"k����T$T4����U��X!-ʵ��v|�*c���,�o�����*yjw��Z���	��n�o(r��l�MbUu
�����h�9�^�dя��#Qژ�4��篸3fw���c0�FV�K�;ǡ���^h1�
�J0ǅ�ӎh���bs�b�� i_u�j��(���By�q0C�9N��B��~���r�#紬AJ�3��$��B籦�ZU�Ӈ���)�$��%S����8cY�%�	4����B\��r�8]c�`���S��H��1Mg��>0��qn�gXv�eP���Ҕ�$�X�)��Y\��K��}����@@�ì��������G}g	T�����3�!��m�qN�x��Ǝu���PtKE���>�f7��ګn�h�i��r4,I�@���1���-03Y�ZdR��
� ��B�� �hN��P��@)�����d!Ø��
|�9�)��X�&�:K�9�=��R�z�,kK����f��b�����qA�{J[غ`��~�^�m�?6��p[�{d/a_�|�2{�p����j+�mDTb�pn�?�[�� h�qw�2�|�?L�1�w��g�Z<��/;�]�4iH�kx�>t�s�D�a��e��xm���խ�*�-�WnI߬%p�u�����ÈP'�t�Q�s���c:,�r�G>��+|[�] �}Ϊ�?��l�ilY���R�X�Lig3N���� �Y
��kK;7|�}����ݝ��j���H���w7T�\�w �Ƀ�J`)ys�a�z�Pp���z�!^`� [?�t���u�|Xz�^���D���\��^���w�>(����f֥Q�����4��u����!�0�����~�_�\<)/��uK
ES����-���j��z��`Z���oDw�r~��T�UՊ��=��ߦ(a��΄kF Oa�J���Cϱ��[���88id��ht(أ��!�}@����qs����Ό�I&ܮ�rI�t���JW$�d���z�S)>E���4E�bG�sB���L7�̮S����Ow,�OP�O  $l{�����&S�8�b��?��]b�j��{G�;�P���*M��l�eC2o=l=�N
 �l[���+�$����:I�0�����2���kւs)��nfl��]YeV"�UZ�$ҍST��\�9�;�{yn��ߥ���߶-���\҉����}Q�	V�Y����ǅz�z8��FLF$�Q]6*h>����>��cvC	[;�̣0pz1M����¢��b^���r��'��".���nK��c�x�':��6���J�`2lR���{�`衷�yS���ͣ�ݑsPV�!{m�.�՗��tw��0:�P�'H�p����i���{� ��5M{��[�3�������Mz�u`S\7pF6�"�0 ���b���Zk�Ï,Z�(ԬG�p���і���r8���v��F|���=�:C��驢q_�!��d��'�3�n��F%�	���W�%����q�|�
(,��D7��5i�c<�+��-�=Y���^�!�	\#�+�^���6��W~�m���h,�1	�rSF����S����^�&*��+�t�����V��;�j��H�&�5�Q)K��r��!���H#A���_֬�w������ �;&��fI�"��k�r���:������R���p����j�����@uT8{�w$�>���UN�d��c�� W�����������l���Z(,���21�@o���XlOno��� �^9e���/eaSm�3m*�=4����TE���}��~�F"�U1	�%�Eتd=��/�pX�(����ru��4��-�x���T�7�]"�JV�r�?ȪG� �ASpqH3d����+�&�w~��&!�\U�M]G����eT�8�'R�߃:ڹ���%8X���1��mD"�'*�+�*��i[^G�����l�xv�Q?ˊD�Dď���A��o�Zc>ju��:��sd	�v��! ���|���K �WNQ;��#�Kh[��(fk�|1k��]1�uQmU��V��a�o7b�ZD�
e��{�3��ԕ�Ubj���L :K~�o�v�jO(/P�!�PԂ˶lL�Q2�x�������.z���`�(�Y�|	0�#�������AX�v�%vKD����̓�[��K9��g�oW�7��v6�GC�ڄ�F�wڪ�#gl�*�7��E ��ٳFdԏ�*�m���	�|`g�S����4,���Q
m��@�g�(�I �.0`�Jy�TY���MWvǰW&��{�I���z�g^�S���?zt���1@��bf��c��>���PH�P���0:Çu0�&~�%��ak*S����tٻ|�u0x���!�\����.�
q �[��D�W���fģ|�o�ti R����l�mqW�^0ku����"�~��"�R[z�KNƷ�S��h�mj�3������a�O��B`R�G� ugn��:�äCÀ�BQ��Ϩ�,�������ۇ�
.8؟�d})�e"�U�Kn��=4B�S�x	F,$:��rZY'\��mav0?�H�ZT����<b�>o�|��WaxF[��`k�P��+���W���WwVKy�uw��B�ڂQ�qm�f�
�Ai3H.G5Cz�N�:����I��ռ��xx;A�H�Z�B k���ld.N���_�
}P�R4������=fi6�FD�rW� �{rk8�j��>�P��.~�/�>̖6L����-�l�6ǩ��#����U��8���q5,����]U���<Dۗ ���Z��.��i��c�9��UY�,���v����5b�yL��Tb�e���d��|!A��O���@71�^��Z�#� �*��᰿у�b�TТS��rS�&��[*�:{�~(�
��Riu@�8�-��T(t���a�-S��^���<1�D�Zl���/���g*�D�����XX�^d�	�L����,�!Co:��c̝ϷVM�O{ {�褚�ث���
G6���a�Yu�_k�2�H`˱���#� ��FI�}�3��� 4��yѕ�(KU��b�o���ˬ�fd��f*}u&�s�3�n�/�Z&�b9P쩪��Z~$�_�3�.]�֩A,��_<rJFQ���@c�e���*��(��N�Ɠ���Iмތ�Б�N��Q��.�Q�w����O�,C��BG�er�P5�l�=�(��L�n-��{����!,�XSA������b�Qᅅ
Nf��a��X��'.��`�.��i���C�p���]�P�f�b-Ӛ��I �	G���J*1���8��$i&>�קU��0Y:�d�����R�7/���{�3��wS�c�;���4䊬[���˄�׏�?nC9�n�`�W1-'@Id<�����Iݼ�K��.h<��:>��%Oç����a�������$���l���f�kx�n���ͼ,�P�i+��=�˟W��\�)nq�CN�ֵ�H�i��%(�2O���?���N���R� ń��H��D �;\�f �kg�g_�a0���Ɓpe�O-r>d��Sְ��|Yy>~��M(�zq�ro�Gr���+N.��Q�=-����@X���VG��U��}J�q��|�o��^g$�K���$����N�O_�
�Q���g�ț�&� �G��	�$/`��9t��mL���O����J]-$�c{L��<�xǦ.���,�fEa*������r$�_2�@2�J"@�C�A��olg�F���D�ً~�]�艍Ι�g]�a�aU�{F� 0y��2h�����%`k�1��;~���CZշ�y��L!��H���C����ZR�.����Z���H���DH]Y�h��%
m�TDɀ��]243;7a�R���/����h��m�r��&��'[~���[�9J�ձ�)4ku�4����aA<�=i�侓O�l�4,�}�� �`��|"��~*��ޞ����!M"�Kn�g�]��o��"��������}�3E�uD��p/oh���1��;�z� ���%	�:�k�x7���Hz��B-��?�m �j$,cIn���rT#�K���L9�K�����H�5H(Pw��J�g��J?�鍤�­���|��̑+ͪ��/��#�V�c�:�Yo���j!^�W�	x�D�hJ��%O������,��I23�=1���6��l}{DW�]G����l����FEf�������=M)���8Ʊ����a��]�Y��ˁ$�:�Tt�/襷N����kɛ�mF���X�&����+��E�(��������Qx55jk����uM9�M��O����/R�@1A� ���Lm�;�$?�k�k(1!:!�%��.r	L�y�R��~W6n����n��1
峅;���01O!J�'a|�63��p9�p��@�AN�1�H��T,$7��q��w)_V�j�ճ&̈����hѧ��G�B��*_ĺyIm����[r�5Z�Ld<K#nLv�إ����gO�N����|[��~��a��#�m�����L�H���8#���`���>�!�č`����\J�