��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����N~@#�k�0!����+��=L���0�ԴZ�2�Mc���ZO�����=�����վ�	"cqw��a��TS[��{=:�����K��-�մ�(��k��N�-� 偙O��QZ��~rL'�x[�i,mׇp���O�I43��4d�,�H�����SN��d���3���r��m���̨T�I;uj2Y� Er�*p�Q$Gm���p�V�`�2^���,hz�<p��l�Bxt�5��s��\yq���#�@W���f:m��T�	,*�񞭋����_��㧋l�	�\�:��uGd��PǷ��N�I��_����Tuv� ���us�(H�~�{2H�:Zor�Q	#%�3ˠ!��iS��95�,?�.���/�F�i{#���Tp5����Ҥ0{%���2vpn���X�����@l����3dc�ק�3	�Ed&3�ZN O���z��s�yxӡt��v*}ԫy nj#��lc��m戭k[��5)�A#�����8�!�]�Z�s�M���t��w�!��'ÒE�rv��Ϝ�c@<U��\tq+��&|�&X1)C�����r�A~��B�&�����s�:n{p��͠R�X⺂L^��R����c���f��J^?��ܣR�O 1�rV���:��T�4���AD����˩�F�w��)Dm�O�b,�a���1$��c��7t[i2>�ޔ0,S���󧇳Ϟ�ᒨ�-��}�!6��Jyv�醊�^_�(�H�(y^����o#����X��3-�k\8�M�T�"`R�DF6ȕ� �,5�;Ҭ C�k���1\������k�t־9�}���� ���QHF��"��t�9 ?��{E_�7��!����](�S��0�q��w�9��=�i]�1�GʦȪc�W�XC�|�$��}q�6����zf(����լml�dz������*�eLD�*�,�m�]ہ6����D�Gw� �g��' A���FX��\өܹ&�6�h�Ð�$�(+��埧��= Eza ��찠pr[�c&��nP��x�2�TK�M�V���3Y4vIR\������ɭ�1՟?4�_y�y+����ƄJMm����@����m�����c�t�����:ud�Q�����T4���QxBŎ��\o���t�*Z�$�*7<�t~eP/`lfhg��6��[nn��#<����n�D:��pI����ߣ��P$|#{�������]��?Q��b�$~a.�r��9��@/��:��K%�DP0�}Pt*�R�1��5/f#���^^
S2��|��L?���v��W:u}�b���,EL�t�-*���{˗����K3!��$0���$o��|FL�?vKƊ,��?+�� !��Y%�F�֠yTE��,�2ثÄg}�L�=v~�2H��G�E��[�"1ػ 9����s���kF;U �f�d���7Vv���FꞋW�1�n�-!LE��z8֬�{�D廚12njp��N��Jg�v�u��J>��:�+�����yB��Ǝ�p^ �=�E
G	�-�Αl�gXы��_Z�g�1ڹ�B*���i���(#�>]04u05H���ӫ�e���C`=|����:��SL�W�]8Wy|˻����ԫ ��_$c��(w�z���{�G��B)xɗ�6��n��n�	�/ܶI<ǳRT=���g��u	ΰ���,��A b��Zð�y�O�#XR�~�RN�شfVd~̍mE�g�;"��F{p� HM�{޻�^O��N������ڎc����,���1��&OPS��6��>N��s���4[P.i�-K�� #��!��3��T]��׆�iч�iy���rE�5�b�)s�Tz߸zO�l�a�_��� $w�+�����!F��xL)��Q}�K�5uhuj�>��](�s_�Am�����'YPqI�M�3��hx;��9{��^p�k���
�$��3B�}���p1���8����9X�(+��R� i�H�Xg�#��Ҏ��e�1�b�� 0)�6�p�ܚބ�� ��a�h��^�M���uXȆQ�b�3���"��:��;�.|��������<~�s�2�W�"0��Y�^�$�S�rT���GeU~���ޛ>�2\��������&����o���B�K���)"�V���&����YO��0�#�Ft�2Yk��w:I�M���ᐿ]8n,j-�P
\�k�V
�~��X5�Ӱ�z��>k��s ��g�1k� g�a�5��*�������?�������4�ӱo3�{v��N �~�ҁ8�H���nF�㥳q��3���t�܄Z��>7*(�X�B�nm ��a5�C�]���숹��W͡��� ��p��� �K g�*t��o='(�rg��`0���N\C*&?\T�٪Bq^�X�$u��է�Y�?W�E�%�<I��y����{�mȌx��W���G�p�;u� �!N.E���+ƿ�����|��g���F�\�&eUx�O�x#=�"%��n�V�)6�Y���_��	L�����D�����af����2�ic���T�:������EP˰�d��tʺ9ڒY��� �..�s��Ij��Ɍ�,�g���57���=`��%<}'�8=<N#�r��У�C��2G��R)���m^s%���|���Ki�E�ȄY�oN��ssY�v�ɜ\�I�[�mB$J�D���U�~�z,��GQr�.��d7��j�P�4���q��7�5uNb�Ogj�	�DU�tE�/{�*.88YZe`�.�*���(�5yy���Ġv���M9my*���o�׌2�u��[�:V߃?�W�Y��3$���K���m��w�5���a��[K��q%	�E7ļ�ԍ��l����@�������X5��[��w�t�`:��Q�3�lH�����h�����/��(
7��I6o��(-Yh�1��.���j+�c.�m��-��1��ր�YM9������ʕ�a�o�M<a���o6/� ����ٳ���F?ra	�b/�0��e�Q	a��	���~�̈́E,g��#H>R@"�[j6�i��!%(��W݁	��%#o#�}o��nV�tf�z���)0E�JQk�ڳ�2rS+��C�f8�;��)�F����Ŝ ��e��<�Õ�@Yw`�����'������TP�:ؓ�vI�_��`���!��ͩ�1C��
n����bD���&_-�D���մ-������d��a��8�̔ � �����V	����7d&�XM^N��_�qU��/U04^ҕ�; ٟ��v��؜��R�ߝ­"�9��D��L�/4��%�
Ȉ����u�k��j��Π�Ư����!��MGA��T7N�#K�G�ꡔ��i��#u�F�F��bÔ_�HӜ�Rėz�pk84eY{i���?x�-��ZY�kD"ƀ R�C3��{-,��e�j�|��(�|�i#*�*�l�O�{a�16 �H%?��t��sB�Q�	k�
8�Y�u۱�MAGN|JԸ0�/GS�Ԏt��芌Ch����aw/9�у[�	�J�p6�w���t��Yf�ߒԂ�H������v@��ĶO��M-[!��0OD�����T�q~*��1�&dG9%aa�������iζ���RܕlkP��\7�3>�d�HL�S;v��~�����Jv��|�YP�<�(w�S3����Q>,�Т哙����AW	��P��FJ|��{