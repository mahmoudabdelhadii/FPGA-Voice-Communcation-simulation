��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����N~@#�k�0!����+��=L���0�ԴZ�2�Mc���ZO�����=�����վ�	"cqw��a��TS[��{=:�����K��-�մ�(��k��N�-� 偙O��QZ��~rL'�x[�i,mׇp���O�I43��4d�,�H�����SN��d���3���r��m���̨T�I;uj2Y� Er�*p�Q$Gm���p�V�`�2^���,hz�<p��l�Bxt�5��s��\yq���#�@W���f:m��T�	,*�񞭋����_��㧋l�	�\�:��uGd��PǷ��N�I��_����Tuv� ���us�(H�~�{2H�:Zor�Q	#%�3ˠ!��iS��95�,?�.���/�F�i{#���Tp5����Ҥ0{%���2vpn���X�����@l����3dc�ק�3	�Ed&3�ZN O���z��s�yxӡt��v*}ԫy nj#��lc��m戭k[��5)�A#�����8�!�]�Z�s�M���t��w�!��'ÒE�rv��Ϝ�c@<U��\tq+��&|�&X1)C�����r�A~��B�&�����s�:n{p��͠R�X⺂L^��R����c���f��J^?��ܣR�O 1�rV���:��T�4���AD����˩�F�w��)Dm�O�b,�a���1$��c��7t[i2>�ޔ0,S���󧇳Ϟ�ᒨ�-��}�!6��Jyv�醊�^_�(�H�(y^����o#����X��3-�k\8�M�T�"`R�DF6ȕ� �,5�;Ҭ C�k���1\������k�t־9�}���� ���QHF��"��t�9 ?��{E_�7��!����](�S��0�q��w�9��=�i]�1�GʦȪc�W�XC�|�$��}q�6����zf(����լml�dz������*�eLD�*�,�m�]ہ6����D�Gw� �g��' A��)�m���b�����L~�B�3A�/15�s�dm�\��rbY�6�g��x��E����Uf��)
^fd���YaŌF�<���^1!�C;4�i�@��e��f��1GY|\0z��Wea��".��������Q��F}zm̋�{�h OSK�&y�À� Q������e��5.��ѬQ��G�P@��S@fx�f��{���A�������U�ǚb]wT�sS��֬���/�B�'����	bk�U��p����"�-m�U.+X��p������J'I�^�6��?MwZ��ݭ��E=Eu'o�#\t�>A��:Xۋ�G�ӎ�B��7�y�4�)�-��I��"�z��̦j��Ș=$ؗ5�%��	(֋�f�\��w�~��	瑡��aW��z������W��P�t��cq�0kXnG�� ��aW�	� %|ꦙ�����k3���_6�Zxsu9j��>���bGN���)��Fߦ�Cr��,/X�a�3ʨC�{��*Ɲ��<S�s���ۻ닎C��I���(�BI�l���8U-��;��*B��ӵ! l/_��?b&�^uN�wM���T�L%�0�/Y�]�q��S�{�E*�B�_b���%-WN��m79�14�D/8��HJ��h�lZ�6������0^�*��'��/��+����� RB��F�5��O�)�<{:��WYb�uJ�!Q�n�r���
9��s�6��c�� A!��t����	:�R�&ҩni;�=�͈���j�`���1Jn�g�[�o�dkE�h+�XX�
�@r1���G���M�az����X:-��Q,eu��湞r�2��?\�~�xn��ڃl����~���/����
(�d�只�xE"ӣU�o$�ol.�{[I/c���E��� �yqe.�3D��� C*����a�C�r��I�ôUi%��H���ڕ���iᕖ�4�n�t��."���",��5n95�0y֭�V�����nD�Bi~H%fyf�b�p�}�~YH�V:c��WW��7�d��W#_&��D=`�f�"&*��],�6�@�<� 2�j/ �T68K@�ߛ�2���i,ToB�}ղ !�j����<���l�ړ]�3K0�(e8�[�����F�̈D�|4����s�(�Ԣ����&�b#���s=&c�X����~_�z�ӷbf�;��H�+,t��ہD�X��֦��"wغ��Hl�2H?vRw�83P��PݙG�GieY��A���Y��q���0vf����\�1�w�q�<�R�9t��~&[?��Hz��Rj:�1�f?}�����;KX��z$���C�\WC~��eG,�_J��K�Jf���ZّZp:1�k,3>Bu6�XwJ�x�w��a����\6�@S�x��/M��x\��Q�&W��WҰ �08ct�+''t���؁]�G�nt䶔�(�;WJ=�IҸD�S@R�VVƘU�e��u	S�p�7����e+���ٝ��g���>R�K9R�6$�c��^��YA�n")�?PB�:�8�h�e��7+�J����x�$���\��#t^������0��:Sw�Qq�<P��0����=�����V�����+ċ'�Y��,"����ۗC�&��Tw�ȕ��~`'��X� �Ia L��M
(c����;9R����[ZV�L�Pg�M�C��~�4�˅9�����ڑ��|�����b����~	��1�,����Q�`v(eP�7�Y�яh(x�Y��s\�o��c��l�`>}��ߋ��Z�K��u��b9*mb����`����>��R�r�-����q���=v�XŲW
�ȡ���+igJ�d�1gj���j��Y�̜��r'���-�����NK��&@�.M�t8�� ���^��/�ZZ��3�r*$���2��8w)���&B�6�)Q�Ҍ�	�d��@���G.����)�g,�,I{42j�B�,{�>��ٽݨ�ܑ�}SD]X�������|-x��N<̒�zz+�XEWR���B�^�@�%��f��]�Vm��wp�����<CBc�T;aO��n$�x6"��}>cѓ)��^ױB�"�j�1Tش'烃�C�w�)�)���W����|�A͝��E$5�~�xv*�}1��T�^��� �C�D�幟�f�U^���7n5َ���S�r �Q�9��(#XmDY��P��*'�6�����r�0Y:J�z%
)+ESNU:ex�kfN�A�*�#��땊�ߔ&�ߋR��Zh���ia��7ӂOuO��X{U��nnm-��`���n\���[�'���u���8�C��:$���/A<��3�����t@jM6򘸝�T-�r��c��t.韰�~� ]C��|��֓ں) �^p�]��(��%"������,#^]�s����}0C�bTۗ7�t3 ��d���p	�(C%e�q��m�x#������n@�7�uN��F�+�`H�h`��,�.9�(�����\���<��u��t%8�z[-��O?�U��<�Ѝ�?|�0����'��~�w��9�x���/K��{%շہ�J��X ��C�ݨ� e��%#��~�?�����[!/N?�ޫ��K���(��)e.�h^�Vuw�4e򱨲H��h�LBJRI�a*��L��5$nȾG��Ӹ�LD(���'mP�u.랴�2+��TI��_fݠ��Ѻvi#n�? )��_
�T��A裤��Ӆ��x���@]�
T����~ 6KO䀐�"3[��*�	�3��Z�(� �ː��m_pS0v���#�')�B��_˦"|%�tp��U����{r�q��q\����N�Y{H��~+~��+J�;�
���l�ڃ�ۡ�eZ�@ߠU eT����"��~7hk�+{L�Pg:��E�_%W�ջ��=N�)���i�n�<m ,T�E��c���\�����S����ʮSH��0����D��VD�룈�dQ�w�M�q���2�+>�ֶ����ꊲh��(�{y0�����f�w�r��K&��� �[u�JDl	XI3dB�^��Ї��s���'���F7*��F.���7��5,?��ژ>�Y;�>SNr<�!o�5�>�����9���~Q�91 L-��/��+՚(�틷gx�5gP��TX�0�y'~W����R�c4<%;a�mP�Of	_K{�2�"�X��ž������ʽ���Kwx�]��/���'����lP@��W~,q�맿y|3��a�|�6�|_z���rk�e�;�P4k�t���y�?7����1g:�Hˊ�.Jᾤ��M�����X�!�ˍ%ZwY@T��-��^J�����	�~aT���x��%i{��J�?N�Z.�_g�֝QB=���~t��{Q-E]��fz�,v(-�t]sE�0��esu1.�4�����!���:���IX�1&C|�T�/�l��9O���'F�Lcކ�&Կ��z�;Pf+��%��@I�ћ^3@�ämc���g�*�ۜ���9˭�������.<�*B*l�R>,�M���1�	l�BH�8����i�&4�N>v�"W�q4�;m74���1	 �*�7���7��g�#7_�^|���tϔ�8�9�f�~dT)A'�����ULA=�E�h�M��Ϗ��G��s$8�q���CJNͽ9P�%`9q����,�+j]����_|�є�uEñ7uA*��:�9�8ޞ�)���z;bls���ydO�<����σ��d��N���߭�z>�ǎ,�~i��l۠��"/���m���M�S({;����?��1̍,ra���� ��D������j[̍�>2Aǧ�O�zi�$��+3�-$��<��r��-&�04P̨|��+�����H��>�a� �����nt�|��#xn���D�
VU�\f�qy�ՠ,���H�E
B&�s��I� ��Bs���2�)��Y��-�%��w1H��E~�