��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����N~@#�k�0!����+��=L���0�ԴZ�2�Mc���ZO�����=�����վ�	"cqw��a��TS[��{=:�����K��-�մ�(��k��N�-� 偙O��QZ��~rL'�x[�i,mׇp���O�I43��4d�,�H�����SN��d���3���r��m���̨T�I;uj2Y� Er�*p�Q$Gm���p�V�`�2^���,hz�<p��l�Bxt�5��s��\yq���#�@W���f:m��T�	,*�񞭋����_��㧋l�	�\�:��uGd��PǷ��N�I��_����Tuv� ���us�(H�~�{2H�:Zor�Q	#%�3ˠ!��iS��95�,?�.���/�F�i{#���Tp5����Ҥ0{%���2vpn���X�����@l����3dc�ק�3	�Ed&3�ZN O���z��s�yxӡt��v*}ԫy nj#��lc��m戭k[��5)�A#�����8�!�]�Z�s�M���t��w�!��'ÒE�rv��Ϝ�c@<U��\tq+��&|�&X1)C�����r�A~��B�&�����s�:n{p��͠R�X⺂L^��R����c���f��J^?��ܣR�O 1�rV���:��T�4���AD����˩�F�w��)Dm�O�b,�a���1$��c��7t[i2>�ޔ0,S���󧇳Ϟ�ᒨ�-��}�!6��Jyv�醊�^_�(�H�(y^����o#����X��3-�k\8�M�T�"`R�DF6ȕ� �,5�;Ҭ C�k���1\������k�t־9�}���� ���QHF��"��t�9 ?��{E_�7��!����](�S��0�q��w�9��=�i]�1�GʦȪc�W�XC�|�$��}q�6����zf(����լml�dz������*�eLD�*�,�m�]ہ6����D�Gw� �g��' A��)�m���b�����L~�B�3A�/15�s�dm�\��rbY�6�g��x��E����Uf��)
^fd���YaŌF�<����^ڍ�-�L�A�hm�Z���JA�&�拏Ӻ�*�=�#��Po��[U�Ƞ���>�-:NM�)��Μ&�^[\c�s�.��i�����+�G'Y�h�8�|��d�j�?v�,�e�Qy6p#��w%�J������q�O�U�>�(zHO�r%�`V<�Q�O�+�Y"��9���1����zlP�
�#�i7`Vq
|F�L�-��x w�lP�)KG�m1�V�Zq�����"������kjk��8Ľ�h�akF��� ��� +���m}�k��r5%�k�(yW1��|
}$�AE���s#s+p�s+F�����G�1�t�+Q ��AO� e/�%�k&�6�t<�"Ln�����Ps�'~<����h���Wl��]݁��h���\�����62]��V,|,��W�`(���ӽQ�.I'���#�ez"�k��F��8F�H
�P���u��ߟ5�*ѹV�x q�]K��I�X��xL��4U��i1�!�
H��Q#Z�%�����#]�� ��dV�@�6;9`�+Q���H�'.N�c�������K
s�{BbJ5�	k>��e�a�6�c#�8�C��r�9gW��P݆�1��¬!���k��6�]O�Ѥ�n��t�q�gfK���u׭,�S9_�DB�x�����\���qC'y���*�/s�+�(*_�hR`�4������EYt#z*g�9w�Z举�s?���Z��]�a�Ky������{���h5^������^G�Rj�D����A��N5|R��K]�ջɬlo>8ɧ>�)9��{h��c�ҟ����% {A��&Nʞ��m�b�2�V�t}D���q5�s"��dIS�m+�?���ɬ���_(U����MMj�WS� \h�v�W�J��R,L#䬓"
��W��8�ƣ�L	�z��c`�!F���N��Jr��4/5��-��G�ܧ�(�x���}�cw)�R�����Ԛ��SZN0��6��Hxr}�Ld(o Jz��[��L��W�C���>���ZC��m�Z[��-wW�g���10��']Xkn6h��O�/��H�8�Y�`�_���S�����z7@%WRr��]�Y��%&����!i���&���R�H��-F���h��T�0��m�2����#B߸����I��0�S�4_�A!���E�xǚ׊���9����F���
 K��r?	��d��5)A,���J�.�ɖ/����]��sC�l�d��F5��<�tS��R2��ͽ;��������0vu�_�WI�)%�Q��0�B�u�0l�ࢠ��E-2�>^�u��I�Z����;=�'�^�qu�_�y��&D)��g�Q1^��i�(�=���% |sT��"=l��I���Ս�,	��RS=���[W��������s�R�&�R;bo�4�v�q�띋��+|߫9p��}6��}wܵ_���Ĭ
&I�?�y�
����D"�W���#��<�h�#k���W��ǉ\ƺ����-��&Дk�Pd�ﮥ��w����K\	(��a#I��cN����=K��,c2�k3l5)ђ�t2A{_`�������q7�/�mu��B��R�BYb�Q�_I�v+� /K&+��*����/|X�"H��m(5c����>��``��B!f&��Ѥ��1�����I���6������;���F̀C��?"U�(�w6G��[�(���n���b8�M�K�)�3&u�1C������@����9�L�%������S�W&}������h<<Nzl���g TP*�;�H��w��x����rt��-©)C춪���6�j&��'��7��4��:�nD��h���y��B��i�@��K�CSJ���l���[*�գF�DhAe�EG'�^6��b&����Tb��\o��3�vgx2�q����a���z�TR��7�;�v%_�#cl�[��XoO�"GQğ�L�b0����YE-� HL'1���9ɯ(��O
};�DLjCQR���4��v@T]%�/,� �.���ds�C��"6���඘���Hp㬚VL,r��<��bZ"@��=�Y�Vy~e���&��zdr�z��|-jk�b�WM�?�,��R�	�Ay��u�~УCc�h�{"]����b����(6r6���}��͸�)�������Zsf�§ ��1���D?����iĨTE�l��R�:g� �h�7WS����XZ��.�,&J~O0�R���>ժ��XM���J�%ZI�TJ�İ�~	6�3Y��.��;� o-;��#���
�E�F�,�Y�>� әSC!B4�&�"T�m��FR��Z�Tf�f'T�����,Yu,����]n��
Ķ�&j)ß'�m�4��&NDc���N�C|1GP��Bz��(X�C��E�wM�����7�s�0�1��u�J�AJ�͋�:��)�:���,(Ph��9O!�y��R�`�ؙ��x����r��~����P�M�,v1�:�-��]�%JK/a���=睜���T�4�L�ko�ہ\1h�{L�ڲ�n��ZJj��9�bY��G����
��Z/?�ٶ'�ED�?����߀�����&�I^m�������^�#��c���&+�v���#��Lx���%���}ꀪ�������>��2&�����A�����Y9 ��������?ҳG�U^W���@F�8��ma�ͫ��=d�����,T�V�T9X M���j52,C��>�Nk�z�.c��V T]�P��\���t9�@n8sO��Ĵ�-{�l�p���1x�?���FD�*҇Z%>y��<N���0��I� l�i���Y��.	��H˅�̯?�+R�K?j��{��|���y@���{�e�� ���נ�����ܻ��n@f�:�`\�%�)Ou��^R���9%���"�6�Sk�]��sCIt��[������������a+pG����NQ�滷�?oa��V1���l2M��l���f��G���X}�\���_�u�$�O��0J�'N�8�$�gZ����y��,�mb�3l�g��
�� /ߋk�9I�B��m�I{��G�wS�W>�4b�䧃��b����R<�d��%��ǝF�f�"_v�Z':X�����w�f������v�:�-��#�2��.���҂6v�^������qm��y;�}f�<5���6�1�i��I�����l�]��I`��3S��U�S;�X~m�l�D5�M�&�2�7�z7��N9ZtE��X�臙���sq�;�ksR��>@3��Y=�I%�0�ޗq6�l(�Lo�2Jz9vZ����9*r7��$R�_cFN�1̅n���|X �f���W�ɩ����aA��z)l��4�I��_>�=� �W9 2ך�l��a��6Y%3��A�W�(y�C��oK���<}����g��m���V��Y����1熣�񀒟Klt�_Ԓu�HD��G�X�� �S�#�~�1���ⷻ�f���j1K��|����8<be���&�7��>:zp8PgK��,�ennڏ���C�-��#��oJǉ��̑jz%`�� T��1s�J������b]�4�=�:��S�Y֛��+!B<�?��+�J8���Di
|�C�Q h�$�{�(���F_����>��11َ.Fn8�MC��H
'�#S"�P6�I�d�e����}�H�B�xV#�e�"Oʖj�pg�d{�$�����(�]9�dq֯���e4�p����4���j#q�t���3F��sn	���j|��o�L�Y#vclFh:,rt���� �批�`�WJk�Z~/�.Y��I	�����p�Мi�|��Q��'��m1�C�X�����Dg���3�Kҙ�����,yD�p����a%��;�k�5g&��!�D�@[!�i�N�����F��z�`)��KY��X�ɬy�f^_��������4�c���y'L�a�y>�x���Q 
���V88C���ŭ�Df��߇�/E�a���޺�ތT@و=/F�`�3��1S.j:7`0g�Z��f��|�
�f��f�0|waT�ʿ`~k�Q�HE��!����9�j���S�)=�Z�*X91��  ����?CL�=��JO�J��~0�
>��Jk�N3�Y�5�����t|�z�-��S��?ʳR�sA�4ʞf��	.�il ��P�>�)�;Z:Q��*L��A�ڛߟ���j�n5u����|��T��]|�>s��㼡�!����%����_y�ϯk"R����>�C8��bl���{����һ�BlO�@LJ: ��V;9w��h��E�����%"HV	o*��WZa�-�Va�����r���S�}�!�ӱ��yA�ͮIIg�E������0�,��T1�K������p�Xkd-�Ka]�����Û4<�,�5s�/��<3�V��qQ+f�{S�Oz0e�U�l̥_!@�b�>�	�����pih���3�<:8�Z��o�+os�w[3�$�i��+H�RL1�HK�Iܦ�%'���J��9=�^���Nw�����8�ōNw���ɘ��V�B��kb1�ܑ��!���!`���3���)]��8#d��Æ�	#u�=�$i{�
Nc1�&��n�*:�gS4��o׀���a��R�%���#U|�t�m�M=���ӷ�[��7�$�!��sV�C��?9-2/@?x�����g�P8��q��l=���x������Z6"ө�kZ5a�:�{��F�@�?"|w{�3���l��wèʥ���^����ȶ�q��6nm�Zmr�$�����x���!#C|��Ϳ�ެP����bݣ�Uߘ�	�!`�N\
���X�
�d�{��|2���#ko�����k:�g���BѴ������#A����h��UF����ئ�G�Ib^��Y3s�D6�s蔌Be��2���Y	b�gLJ�>$�Yu=�!�ܬ�E#$�k:@��Լ�UA��G%��!����0am��6j�Ų�̊&�Ӝ:D�b�]ݻqA��ќm/�|���8��Q	�B}�W$��L���z�+?֣�͗*��lJ?�N��d�x �����F�>�>�˵%и�k��5yi򇭭�[a��r;��Z��;�`	ˏg�A��U�
�V�9=�nTm�i����,����q�!��Yx3���nfy�g�t��ӈ�q,��͇h M]�Rt}��pt�W��7�\2e�1ƅZ�#����w�I����!gt�uٳi5�32���Åb�-�7!��$'t��M��ezuSZ�2Jj�rD�H<r�HgQ���>kK������9^�`<7N�@ H�3�ԋ"
Y��A+�`�6�J?~[F���\ҽ���) })W>t�����䌼ڨf��wJ��Y��X6Q�P��e���W-�/�kx,N���7�����@�ct�n�M�c��a~�c�q����	
C��9)�F�N�AQ=tD���mh�q&�f�@���S��	���9=W��Q��p��}g�F�>�^��[�F@��������3����(���ش�T.�3TL9�|�o��v�ե��g��p�^߫��nӠA�yg?���L��Ϡ"��x���R�z�!��U����A�S�Q�s��`#��=���t%<ʶ(/sD�)A�rn4d�f��I�^Q�e��Gugv��k�۠ 
�f�2�;���f�͛������,"�߿��?��������2���M�X������,Q�՘����S<�"H��2w�I�.��S���-Y�ͩ���H恍�!���7������N�~��uИ���M<n-[Ӿ�/����Vp���ʽǶ����a:� �\���=����I�m~IL�`�=X*��$�a��Y�q�)�;WN�R(&ƹ�J�=|�@- J4�$=�}%�V��mT�c�ޘ󺈱�{&����4������ޒKf#��a�S�r,�
��r�@�?JB�U�h��b�A2��]�y6{t�p�\�]���wW�o$$�iQ<x�+r�ˣX��'_�_��m�b��~K���~�1��mU�����m�w��;�������D��yj8�����"R.��|�<sN��r�<�X��D��������qT򽛾z��'*�#W�o�%��s���o�ӊ���z���/V7���s���əP��E!�uS�
e�m��s���G#<WX���?��ܘ�KV�C����kD1�"
���b<g��^���e��H�mj�cH�֓Kp7�NϢ��e������=��ҏk�&�1V�G�Q��4�HЫOUE�o������W� @m�А@8὎���oP�QL�,�r�b�n��{Ek��1D�΂�c���n�d�(�#�_�<ūE_"��}]������wF��q�?I�.�mm��Q'4UL{M��)��00��H����h�����u��#&�2M���΃������%��Q��Q8x��ꊸ����r��7��z�}fXG�wk��,� PЪ�jS� ֐���+>S#3�]S�)���᯹����'�|*�_���kxO�]|5#@�I�?u<�����A����������1���Hh���A�Ա��E����B����������x��X�K~����P�uu�'S�驗|��wC�ͺesKh2����/^�0�Ł��~�����|�M��E�O�a��p��,�{�Gu���:���ۮ��/v:�O\;|��$ئ5�S�)H����:�D(5xC��Z�v��ǻP�v�+ߏQ�k�S���K�+Z ���k�O!�~����Qy�K@m��H������W��WPO"lIb[|mw�;|���/�u��A$.+*/6�e��o��8�YR����������퓉��~@Hv+93��9c����[�m��7T�������K��3lg��I��0H�l�ѥ��.���"��J�e�U���|�L,t��/�4�_�fO�x�P\�?��'-)�'�c1�ҾuY��	?'g���9"Qu�P�c��,-���	㴃Q���f6FӶ�Hr���4�+���j,�Ų�$nu6\峱�-']��dnw��ʹ�+�~�yER�u�����﬐ZUi����Y<�t0��M}�LvxU��&�uP�v+�>�EJ��_[����D���q�n��Kף~�+)���ں~+Z0�5�����N�SGk�ԟ�$x�:\
��P��E*I��P�Q(�^T\���طD�A"Ij��(M�(n�-F_�C�Ko��ވ�A
�ž�,q�_L uoGT�猍�7�o°k��z>���)?=�a�S��Ӧ3-���!$^�C���B���y����ʴ%��"� JlOq Љ{�8D���͛aDP��e0[���0�J�m����v��Q��s>�G�_�{j�U���̃i�����ڥ�<@�����o��f7?<HM�Ң��CxCNW�����3Ss��p�ѕ�f�QmD���?��vQ.��W�FQͷ�l�&�"�F+��%@X�����F�����}�#�&�]}v��E�Hrr�e���R�hj@^U�𩡩�!�l_�|���1���0�4h�_$��QG'��4y"Q�n�葺��H�X��̱6E��Ľ�ι,��U�:�)�G��2��{r�?R�T�QԴ�2kf���T\t7 ϓ��rX)��_�O��j�&i����n������'�ZB�׎�L��.��" Ϣ�c��R|D55Ufb�_�w����aIk���S�xk��L(���<H� U�T�PD^�e��N4�ƶ�g�I��:���S_�K����Z��H�τQ�>c7W��:p���I�9ݝM�r���肷~��m��CbZh�Jz {b�e���0ޟ�X��9��19)��|_]ʿ��i�1ݨr/����Lm�T�]P��]���j��MF}q�������Ko�.?����Т��#��w(ps�`Zi�L��q� B�����[ϸ"��9��\�_�#��x����p��L7N���I�/{��q�L7ͣBr6hd��JC6&�Sd�ٹ�1��h���)C_�����}��s�f�d��iJ� ��Xg�¯B��?!苒�8W��^9��W�M,e�DCV�vy���Ҋ�������w�=�%�k�D��SYZ���%�W�J@��ƨ��(������ɾ���I�Enp��6��� ��S�K�_[`<"�a�am�y�����(��^�|�Ųo�`�=[�'h���\�v�־VHjv�b���"�.L�"�]Sl�s�qދ]��@:g�O�����~��b�?|�Ac��	f*ta*��"�.CȋmУ@����zY��`wk"��ȵ:;���L_b˪`�6(�z�z��O��5�F"_�S�u���jR��/VJwo�_�B)��Q+
��������`�;��-Hs:WY
���9�x�l��|�t�{���=�.��n��W"�G@5���W��I�@dȃ|��$?:dr���@ˢg>u�j$�g�g�9�Y��B���N�ı�%���`�<�v���8�=٫q�tr˗��I�����\u�b�@T���}���R��,Ygb����R�?9�-^0b��qXiB�[��� ��A_{(]���L���ᤰ��lBb�)�j�X'�jߩE���IC����%u�։{�s��q�$��"[^��%�b�����I��+t��[|!��+H3ZS��zz{��[m�f�˶�����<�L��_�8��lOڒ�7f(/�b�`r޳V�Ý�U,/B��9ܹ�MX�*[T=@ˊ���w�d�y�s׸+��R�
�h�;���0T�&��0+H�f�i�(��D����h�]2�O�0۴V{��Jm�2]R�Ӌ �^���D�V�]Jv�v�RY���๏�M򘮺+b� ,A7�%��|(!!�E^T��YX�9{��� "�Nᘄ3���c6�@=��Y�z ����Y��ጘ�;~��Sa�2��o�g������Q����m�K��y�4ܳ�yz��,����F]�tͳ���R��O#�������H_��5�==�KnS������M�_p"����Y]d�Gn���K1{��iA;��v9H�\�gV���>rH�k��Y>�����H)�g�|��}���,`@����}�����j�^ٳ��g���i6�5
O�ј%�([GE���@���÷��O��r�D���vK�+�ñ����|��Ì�^���x���߳�فێ�7�B�\O>m�y9t��%1.�C����]��Wĵ�q����	�P�i����i����w-���H���k�cj��K!���~^�	�>��-���j���A�z��*���2%W쭱ژB'%ѐ=J&LC�	�=���y� �爉�`ڌ���+�\�6p����Ļ3�&O�>�F��/�ׯs-b��3��85� Vr���Xxk�t�����9f'��K��P�,\�w sf�*q��oy\f��ı���r ��/���$��p ߘ�����?ٵ�Xk�쭅�[ ^9��������=��z�}n � �o�A'VUG޳yb�6O�uنR��1���>�b�w�u�Pj2��P�'��iR���@*�od�O���J0��=G-����P ��t�k�=Y
~�S�FfL	|{��nz�����@g[��i�L�GX���5��/�����V�v�4!خ��ȘL��z�S3z�S�x铷��OD
��@�u|�Q��c�v򼿭I)λc��w��6�Ϻ{�S��i�n}�9��:�;�/;U���N� b)�(O��Q�i`lP����> <S�2󔬐"G�����,���ڞx"�S��]�V-���k��{m�]��ىL���/m挄T�7gǁ��D�.=�r���`�5�g� �9&���34�軅f!��YȀׄ����b���
PHpT���0�̕0	�\�1jg�8���˲�i)��%J?.K���/�R�X�h�� ��XAu��B��k�HjY|&�=��%[[������"�6�E��	��W;'CIb�)b\՘�(�ja�D �����V�q��2T���\X�>Z�{N�8=��xFj�A���+�gx��!L&�I��A��9	B���Y��%��q5h�����z�x��jK���%͢�;���ח��|�N<�,`a�'�@Ï�Ψ��kL��z��~Bi`t$P�ѷT��k��Z��	
1��q�fe��.��i6Ni��J���K2q&(=ؔ�e8��H���
G*��c6~�!�e"��U�m�A�ȗ�F@��eR�)d_͠2sRP��cWĎ��:
�+�]�y�/\M��f�F&'V�+���L�i�O�iP\2�YKF��s7 !���x�������/��lF^��ӉO�q�Z��L���ۧ��eo�|F�u���뿓M�X��;M���㱟���ǬE�
��ڏ�c��~��J 5�?|�V��9��y��fLD���KPB�LP���%V���sp�iŵ��~j6�o��M�F<��%Q���� �h]c�����mͱ��c� �,�#;�9�E:_���t#W��Ӕʿ���B��:��5���0���1ߨ`��Wrw�f<�,���-	H��:'&�̊�����w��@x�)_�D>��m���-<�d�B��}Uc!R�iP�0[<	5�c�.����4
�3�LP/� ~L���U6��H�����.���&�K�T=Y�����o���}׷e0<����<���@~fn0���j��b�^8����u>�@��l[&�Dc��t<$쾚%V|GP�����A�E:)���;�CU$)"�)�Zȧ{�λ�^�`H��6P�&]�a��Hȸt��@C���s� z{�A�ή���z�q���Ww�,��2�E�E��]h�y6��+�3wF��ɨ�\�J_�C_�K�~�WV�	�z�1J�E����4Ж�f�}5=��]�E�ԭ]jw���>�R���9�Ë�3Xtٳ�M�k��ؑ�0���2U���wET�i��h�+Pk��s�s*�ox� ��<+i���q�ff?%��Į�p�9���3��d5ߗ� ����c2"A(�p���.�G���G\� ��М5KgK�_���*Y���dy�?��,����G�0�����ub�D5TC|������c��2<"�=�p��y�}'�te�£,�e˼Vp���܂Q��n![3�Pl���]�]�O�,��1i��