-- (C) 2001-2016 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
rt2U9g1oaqVqRqyVTmqAb7lV3hmrJ6A/qNjbGzDwVmQsFDciBDT4OjEjgwulV7O4LVSYfJx4hqxb
r9UwyaATDSJkyrvxX/kwneDKt/OyzOQ7D6a8w2aKK8QO2yXB/kGpGgykgbsj+MkQN/tztsIgFd4h
dxlTJfbWH5stlxVPNpar0oEnBvK8iE3U8iavjks3q77qIbycZILizGqKhcwTtnyaDuGWPmQbZ3XF
Dn+k5XMI0aH6bAO/vg/d/4ys6xOApEsBi+SjW0ACpmUuivqmLdadnbPiMef/2EboQvmSBSQ03iEv
J82WJ4uEeaq+mLUqZ2qneYdEuaS6ReGFNZRT2Q==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 8992)
`protect data_block
VRwOTX/SfnCxlrj1BIJJqAgOLirIL51PcZ/V2uhZn6mVUtzwUjpGbtAEO8Qlg4SvAXVpM17AVSpC
K90ha55/GrlW9lSgq+/3pDMrQ3k/KV6RozrmPSgRYf8/9yxfsOTxdIJODdFTBFh12TQe7/6im2wI
6ceLtyUEAQ3FD9EZKELsEYWk9iivf6YnXOHKFOD8OeJU/esgEs/TGSqtBafdofp95GgsBmEaDXiY
QCmklUbrDINgk4nj+ZLjIM2tTMaqjkdXmno22RvTxk3anWG5gIimrFIY2A9riqb+oA4qBj+3qd5T
v251mT/2b5FBLMMPCrUsXJ7RhXeber9qAWGERmE3w3OjfL5Mo4+LzEzQL6y+I9AMhOQRQp+f2uJQ
JicOA0RiAKj0DZmkaoWq+BsT71cq9mqFtrGza+N0+OL6l2qB1cAQq4fUNTZrS28ayFXmaYAwXHFu
xxDKhhp/OSfiQa/hEOwEMj3KJ+gTtuiIOktT5njh+H8FkcVGtHyIArcaxn5or871GJG94ZciMfgR
fLzyYvhfwo7wm8IMSqkRUmZ8yfpoUlnStThtkEgEFQBYx6vKRaf2OLjXW8jByOWlux4aqvc3NrpJ
ddvs3ymZp0C/lUjVgNDZct71usLkjg/S9h5VF1n97k00TvBkxXhDbzz3XT4P0ll50PdiyaHtZGdd
XPia8yPp+QcB269au8OdLQMslrWZTCJz//JjmSKV1xNWLySLXHRJc7zi7YghsFFIwCwCZ1Ki6t/7
kCmsA1Gtpo+gOsydOX5CiKjO7F5dIiEV7AXVImiGT0cRsSLtYXqwq+sZB5fOVUsFx462SowkJHO7
GLP1XmQbHhNzyaRPYHm8gG7Fm+at1GshVIzRJEylXyHUOVoXLw7+TfYynf96etc+KKjSVN7vxrYu
3I6Pu/Vrv4n5cvU9YDw0q/RfcTZtzlop8RFRfWcbtJJ3Fln/J9ll7qCklhYktSBquRe4H57NqcDh
WQihU43T+3ZOddRnafDaIxruP2smOjMEErKPYK7WuPcYvlva8FdjGHQoygD8fP/8EQUsyEPIdLah
CAcfVvIIq4HenaH5VRzKw8HDnLcxDNvTo1bImekx3eRQhE7pNB5FZ13gP6Y9ALyvyKa/kxKMD6b+
z9GDY/KpmerJLrEhG7/sS2M7nHtNDiJMCwHw0lOzLZpD8D9EUtVZHOZ7TSx0RcVqwqYOOMTOS/gp
coJXGbjljPmO3zFQgFw9DKPB05NIPCs7sJvjUK6uWOa6ffUT71I16DVIK8Xg306BxCQ3DiNbT2xs
MmBEBEZV6Unwo9x5FuZOxU3KnD7nZortio8gEyFvGhOLPPLCgxfC9CnAIWW/5xRdfnbSjohU42UZ
WA0kV220PPKe6TiI/VlvyqHt4sedxgzvzkXhKCk6t15KwQoFFSbufylCllGItmEZirkdgX5Tq8nv
N+e8DqpeEN8zAp3AFg1Fpdr0I4CsOdRAocWfe/kRx8rgNVReds5R0ii+KcLPSZZDY46nyowT08E6
I5/m4NLhBN1lzdQmJKVkHAryK86kcGPPiK++Ixe7myG/1u71orijGdQ+CpgDZRow2KHJare4+gaH
BIk8aadjixVHkJDlWP0zhelBLAn4zqzJozfbPiLHkMGHJ6amyTwpPBk1U0U+SmnnohTonR73R5S9
TiRXRl0dIYImCZWck4mWaZGvy7wxkMFQ8PMr8c9n5gJzKo5LU1D9HBVRIAyM0ZNyOAMoVkGoL7el
MTh7u1gTQxQkZdvW8skEl3V2b74tpZ8I/TDT9Tb9pkXRw0jjhRvfrQL8ZzYmOyVejADftAwD3miR
xNNtQL4Hr5Zqbo3gTDnb0yvzpsst6w1ruMUqGtTykyNs4KjWxdTFie7WCODdEDzyVhvVImQl4ESy
Al/eyvjw7TxzXEtGANJsv6R2TO1OJBUmKTlFQRWliZeJEIz2fh/ug3fRJn1nqqGqXucwn2hguBjz
AfRFDbhqzwKkUBW6EUca1Bo0bOxt5F/GoKTdvwXSK7Rfc20kodrobt78MJUJz1gxZcD5EoBBr6xb
WqjvbpWfMyv+jTc3Oy4Y8dsJbBqQy+azkOAWPDN2HWg4ciY5SBIKNyQtvguulAuSQ/sha9UKPayR
jEmyPmpi1vk/URAQJJSFuuEiZhyQHrNnBdMXGHvgO79kAtgKhuOVaBE+rTpEEWV+LixfruzQGywE
dqXROvtSVpCnUgZtiPZ1WWxOl0TBJ0ONRVW8lGRe+ZGkONgq8euLGEuvCsfdJOBZS2Tjt2byLHN+
7FlxK3EgVcHuxerhm4kHS6PHhqELWVETDUDqBpvMe9c5VZM5QhdegNAEgy23D1zeGjdSei7FfAr1
0Y6B8eHW9c6V7mlWF/ug/bKRvNuKLJwdB7aqqnfNFPAf01/K/9HQISX47U3w+K3toJCCF/BfDwl5
VFi0yUOpqMyJc1DsD+Je5uY4+mXT5XZZw/70JwfY4DpUD4SqFko4EkcuzBw3qkUihUdz1FH+5ew8
gxuE9zIJowMIPSx3LStwTfb0V+/cEnDvOXS9bzTrc4gtmHtpKnCKy4Gh8Cuv3DO8rW/jn1NxwwWR
pYZ0DrUC2kHB3T7SZeVI9y12r2fkOJEn476n8A7HpEs6XuDOjmDIwbJcUbb9BEphuD9girROYDiC
aMWLTwTSGib7ojrfElyu0J1OMNjwACUQBOB9xIuig8Nm1B7pqp9YEEnc8kocJOw/oqrOSCHNCO5x
qelNsZj/6351qtE7zE1piCOGWQy0JrDDww1YGraAlh7gK5ZlRyMJ48AyiKIUKZ/x2vgFrOmNLEPt
RbKPWKJtt/z0FCCRdNu+K78iqclS+o0i+tIZ4RmK2++0Gn2QPr2cgbMqy/CLm7S+DA7jS/lSS7CM
4YFQhfQmrQ2zeurArbU/QRO3h/bun0OFbzjGGV4uuvaXon2Z8VthznhQPmyhrBACScZ6wGZNmZGM
mNHwmOjfxw/enNzXU+WEOvU4bielZ2O7W31lawALO03Z+D3xN461wB7yN3ut4owiYOEViP7SGvMU
OLCi1eExNuTH6C6SIUrOu8r49j1wtMIep0uhTv9H0jePxwqY3kc+7K7PSXwu/Auj+xbhtCNqIBZ9
9SCyi/SuEma1pPkhvKYfNS483NdgDhrte9wfvk69l51glshEzkeEqq8uvjoFhhDaYoQ+n3caESnd
EpvtQJ3ancN3Es1NhS+lPxrCnclNOj0wmdyzyBSO+gc49oRFTFqmLUmqM88iJEy8wWDqogfcwSkl
41dtW//NXfeOuCOk1Pb6A6uikFV4OCSA0RHkKiN1DkLHwwunqQua9CutX1EFwCsnhg61EU9S1j4T
o6Gt14wcDUbQVK7vuHbrC6LppGsueq5tV138BmgNEomeXuCYmAuAYA7THivTgSP5BMgPBBeziql+
J/wYLVXXpcxuLaWEnFbMYtsXjkdZNLhoI1tdtX8MnnRPF7Ff2gZwyzfxr260DMO+w/TwgmNyCJih
mbpzmB0jSDwnbVaHHjgMr0ZTUs2V7xRnSc8HOIaQqtmCC1x+r+wHtUaQd2s5+N7u64yQjksad4kS
+9DDJEAbiqOkyoz7AmsZA8n9z2VIeLQW2Ep2U5o0OmuxTroak9bc/Dm2BEUeEmUGtjm49ygscEP0
eTL0vrUmLdElat58I5ZbP+e8osV8wMx+68fs4VmqWhbPp9Mdgr9j/kz/7y5Flm8kgrcge/hEz0or
/wVIEDCSkp8SIOJS9BfONv+UOJFHZC64d3lb1iwNuNJZYOe4wnhmDM9QhbqyXhOmZHtfu3R9KkpP
myecSU4plpH70cxX8qmBvZ4K4TTDa/qjTlG5sOduDBwMmTXtG3yHeFBC0+VkLfFHVqEZTm2lgAz8
cPnhrdWtL++SnnaOQzsn7FmjzVm0RujYGK47UpydEEz0+Bf5jWjg5YzWFKSzvFxmjCCkOGwf54yk
nRLQ3R88ZTh+qxFSfFiCHS2/e7UWYko8WQUAugzh2QVrmTj9BFDWgWBUAJa6FzWUDgRPOH8e8cBS
kW4k09r1Hi6PWmhwa/hkVBZozGo50jEG3m7caV/paZXS9Jn4FKtzRR0Y9jYzYsKW4vzdMeRscctY
2J/unggOUiu00XbXwcUgOLG4ZSqOnHt4rEp1i05Z3RlJjjAa/dc7YBRmD8hT9uVGWBbx3RQgNssp
iSSNe533PVL9BqH1PyVPkjvC1g177sl9o47qv3fL7Y1vWK+4Lq8jhdTFZ+zc7RET6Wy0LaJwUaoJ
xAKNZeyVCRwTkftcgZJe4A9ffDtKKvTmLpok6qgYM79/27El1p5IUB13asqYwraqI510YPM4GNos
Yvz7e5H9fXM2snNj0wniCdIoUQaV7W4ebMqKIxlLRfHmedIK8jwsLqhqxJ0sG+UNF9GOXZbX+XGc
UCtuCXyEWpTeU/YuBcjLBHZLKnHffJBBU4T6UEn+SdclQvSmbqO+rBF00fsgTHIN4Y4j/clCTArZ
hS7KlYQ6+c1dJ3yO1fF8o8C/ep/vYhQtLI/LU9LVvRPemMuKtVF4j/6fPyYbTNFI7pfi8fT1GjCw
ItK7b/txFiiZw2qbcwU8r1kZZL+RdoAcF3nNOXb+s/kDKHScdhTtG6VoDMeeRenMLihbs9LwiaXA
iqEPZhpRucMBZw+Ed8tZXtndYpb7qv1r3+XrdUtxmfkAM90RhlrxiTMdaqKm6uGg24pYCOxCJPcg
N67erlns2htiYxVsZNfr4M+KWVmuRnxIyKwXc5DhkJ2DcQiMtYNsj290Sk/aads0hQ7oD2oOj92e
4JPuk0xlWZHakq3v5AEGtuFAy/lag9TOgWLAR2OJQ+Y1P+z3bJW5d7cY2jYRd5Wgx8d8Y7NaYHHd
3Vg508sHIzZlcxSsG7MZ93iG7gazos2qvidDBfc36WkH6IzuyiWDgbAxrqyg+BYELXQ09jMCn99l
6z42GIgh9TypVUrCWhOQxsYzIRQiwN4MKcyhI/duEZyoaQyJQxuwVG++STODac81zvMT9R00OuYh
ChttYEWmMQaC9oraIH1SDQIa1q3Qk4djA5dIjGy/LhXXMMsVJhFACreq6ihKcTslIT1rLYqpkLum
JnUXJ+r75RS/OxQAzo4YFg2byO2WfsAI518+sB/IJI2+wYse2WToIkpMQ8le7B+HHNMAz17+tFOW
cPPCagR5yL8kanBEgpAsxAixc/N+1cwe3/lAHkLhVddDcPUpjqF0fXSFdTAGNK81i+6wcxg1/k6B
W61Rqc/3QFQrcgXZZ2CDFZFtDDa0etSqpIVRwp/zl6hLJXMQRMDKIhQSPZfe4Jy/BitvAAyc2oLM
4p5P0r3d6slphRVqOcLLrPr1g3ABdpcCml8xiOpoEWfyMC/cAatvKMCqErvGdRQ//VxDesVjkm87
oz7Zruf+gq3+10j3f2cVUkSpk88HQr6wSEyVZ1/jApxaM0WNWIejeRx0gx+hZ3N1LTXK6EgOe+tW
sIemz9UMCJ+yXQJ4TKVmtYEh4sJM8cFbMldS98RyHQY/M30crR2uzY1puUeiSpLbEPl0AvbRgwMa
YsBnCPG2Bg+OQT1hr+E830T7OL5DPjWBmA2YR3/YbGHAuNw3BzvAPewwvWuuPCNEVdG8pfJuFztr
nNDo4uPkev1G1Y+dJRR6hRXfIIplcF7GGrxXI7YfEfmb68Sy2T/H3BynBQiuZs/duUvEIMO/aMUK
bXMIVnmi2ScpSiOH+6eh5HSWdm6H+K77MbNcTb50tP33RDBZB/kECNaH9zuiC8j11kN9nTIXBUb2
RIeLQLNtIJ38Fc4A5yoSVOfl2Au6qfMxGOOHSlE+998+7zixx03mP7/9EXr5qQHsBQR0h83BtNvy
GDVVqDYpAbfQTShiG+C3dmp9KTCSzbzRBJc6zDuhu+ZbHF5mFVYOKLcWjGyprjvY+npLJuhtEIJa
s7QL+Ke0zn+QylKQiPz5l4gK3/q+scsA4oW/qQ8nYWi6OlG7amH/SqVV84hg7mNLS+likQ/xOdMi
bSLR/PMpXixjjdzkMeGkS/x8Pmd/iICjI0QNEgVyS3Tqr27rdzdrJVJZ6k9FX0UtD6rFxVm9Ez3j
dZ8NqR73EDae1I9upT9TsFnfXNvYTrWMQB5LJkeojymqogbArtzAOhKjETyqeQNRK4lyqmAZqnlB
T+e4eHAK29ff4Te4IDwkC3aqJWjynesyWmMH7Z4Ga6EfBh8q+L5OrVxf26HpuZYwZ/SaSKRfQZev
/ethyJJ/poZN35kEjX9Is6zZkpEI9VEVrp+VMVdLI1/DruGTZlY4zksq+6GQhtMNXiVEERFG1RpR
NchJOeDcGgfioDjbSwFBf2eWQyMuqb3wl0USWHFGxq5dCHe6idsCKocm2SgmdUed6zkbJ3NZfry2
dph3/Swg6J1NJZYHj/iLSbBtjoERMx+TiFiem93ku0babuvNVzAKpoQV/+LeoNs1lwoSfsNcGZJQ
/H+uMoYIJlGdjhe+IvyDUWEYaoWflkTIPJwnssAoa2RVO4480rKkVWY8Zv09kU8ID5W9dY1LFVZq
TZhBELl6FJGfKBP8GnoUUXnrjXETovqA8xnBYlTML+4esnY9QEUq8fsNyBCH6lPv9F1W5ABamL8E
0bJm/ldaZPep1daQFnEDeGdYKQno7SrHrS+xCko3mxHkPNY8ErgOVSbgvicSCKEs03pBjQL3pA4T
vQjyBKzif4k8JnI0NFOIzOUOrJKrkeATXWDgkVH4yuKNWkEMrb1Qs+Du65e19mCix/KLZ4IhNftt
txxUM7FM2G/xWbURGgRfJ7AyJm9Wlb9csB5BFroWPsfs5jNmrtmFD9nskIMO5pNNgCZ5nZjmkw3E
vptHFHKFSkvZu4Dle1h4jkEkihrCNSIoavbe56eFlhhurFwxSrlY81dH3/jJff9JAgXYEFCyypow
wjvR/hMW2ZJ8bE9ewHo6aFIQl8oDpurycY7/HJdcmRhYcclIFWS0mRsVdE4d5M+PKw8OlqQ/QY+2
f8/0Hz4Y9a+3fonf7itfplI8DZ7oGUqyUrbhxyni/tgx9Wri1lO8oVBWPlHBv4rXjpvQy5yOK93H
TBXzkD2pF1riVOCrR3cwCtDFdwqs2ciq8qb1ddps6GNteVJjJzM3ZOIWa71zh7uJRGKOH7rIBew/
F6NjtEu64P/WDGtkTgOuU1keOlzXVkWZk5B64SIFr6x0XcvIYcxuFpjVjPZtFOlcUVow7pCJn7Bz
d+D2fq7ypROqvUfYcV1t0+uPX59UUbNiV4NbXezYJYXpdv4r1YwMInSLFf2vlJeNt5GJWO+qxfHz
YpHbOTPsrj10n6rRoDN1KC2gIBHNLeF0wD9WlAETwjoBBCw4kvi2rPj90/yCq8q/pzvAzwnHnQrB
o8PD+vecPL2iGsXx9YK0CoEa3zCzoXUA3r64+hKSqdLjMDaq7/4zel5LnJE6m7iMbUJn7lkEbOZQ
KjLBaGbVue3XpsL18spEK9TowOofHb8Eq1T7vkRDTdYYIQTto5Mp4RRTg73sRTj+5xTxCLL14waw
p9xnTzveoAwquxr1q4bCQlSmPn/Rjb8CJ2BKHnHDCY1AiB2zepsttcMB+4aQSHcZPpiOXidFyZUg
j6CkHiX3VyJrSHM3mJE5LN37g9fSOQFOjMnQeEf/uTB2RUepnM0WqB+fYk7oZ5AmhDJvYmLoWVqU
EzvuQTa1fqp5HJVSFkyRbva5026yVM4GFg0JlFCGjcTa1k/icSRqWmcr2J63lmZ5e/aJNz0Xts6M
Ld5rdwDJ+E3hYegRvNYCzgEBVqLCLuWL8rNVU7JYdK3kTAHYmzNw6JnjW5avZ8AJIDAhobaQGBLe
U66VwN6kBbImkHkaCkgtHNNuZL8Dx/izHrl43ishhVMHgy9VNNL5tuhOSZ6OH8u5M+Ib95eBO3LB
b6P0g88tWplK6Mm21xqbbBpULzZHG6V2Xz7YxPRsZEAx2PAMjbX+ykBIGpeQvOabSl2PzZZl3gBq
VUa6SEZUn4DG0UAMbjQd6zIohTzpQTNZif1ll7Kek8ztLM45ilMaaErCytL3u6mFrfkp68nKx97k
iTYwYfCHi3VQ2yAvCfqKAvwUV1R01yEU75pfeZ21ELd2KM20skOWRV5NIV8cAx6R0B8pRQh+8mxR
HaNDosZSGRFTEMdiuPg1IR8yisN4cKKv6DlKpbYNVubNMm6kyPm5f0pOUhQsS7SjBQIUndSN+HpF
7wYfgkPXXREMYzQqt3ZtyhYog1I9B0cEspbKbPM0qj6z3w/U4vz5/OeLVwnHGTHGLMcZR2uef/LF
2HjghVh5WyGKpLRQEx0YVa93MZAVYBcLLehxTcxILchdep/w4AxQ2JIc2zUZbMdoxS3bqSzZHc9t
M37iuggTR9eA9dN8XZYNdkOgwHKn2YgvkftD8oi3gIcqTurt8fVCyDw8Foxg0S+NbNMgoVZsleWu
GtjR7Q3WzKRs/CyS1nJtri8MUS5O0nDcSyJES+3bbdvpJN9YvqIr4JCL71AmMuhnT4x5G7ztC3o5
sj4kokx3ndIHcVVGSoHtmNVYMVusijQV+eIhlIKgQEDtN58yz1WUB3Ie6rzDWaF2hnlFx8e5sbi5
ZSuNklBrX8tHOtnFB5j4XvTNRonte3eORPtA5e1//Vd2o3Q1q+aaXHmoBL+j9WKE+vjgBlgqfzpz
XVE14HckKmcgPfVc+Tsfl9M8BMBT/GFA5tI8/gPbFMFbOHr9Zny6regPBx21es6HiaKiGjoemK+Y
2GMUBEVIYauo4c4Zmtp9+eHmmV2wGi5qMJh/mIESXt+FdYD1uDB5da0Vk1RbozHVetSKmwec7yiO
FSVMC2sYoxcLLBT5LOcgPit8Mx9R1HvFG3nD/STDdsxDeioZcjdJHYXTtDHtHK0OEFTjFyyMiWz1
AOFnRcGFjk8oRHhtlKeWIXTP9mweFOnPmkmy96RGWCAZk7be5rJo+OSEUJZAfxk2iR7e6tuSmqEO
P3bp0qW1H5Ih4KQUuIx4n/zwr9uIuHCf5qTPBdRDzF0/sM7/ClEw5A3APMm46x7SXR3YO64NUlVz
eYjDNGvzB89XQWEasjLQVvctdUu33uwsHvDK1V72m/jP1UoswRn3Ckkzm11HRlR3S4MpJhdJ69TX
vF+0FzJgykZbtL4HUoAyVhJdQo+LTTTWANxe8u4q/jI6f3QhzBBlC18EFt9vVm2RH23lxdjt0285
dSQdrfGxezaeMlzRadvxFhRvcBYL+jXTl0AuTTC1Hy8sh6EIXD8O76cwTXP82HbnehSW6JxgTxS5
04CJ/f/v5cfzoREzt+BEx9X9YwiwxLKEbizj/9rxWC/HLiJ+rvJjrchzIldOf3ND0C17R0UAZ7xW
4eUCKy6H0C85rVi2PdMh45fu25TMUGhw9L02L4o9KY75xsP031yE6kWmN4vUPCfur19uRgVlWLG6
gu9bCrE0OtOSnRsKMkIyUerif3gsNqVrcgn73KNW8ed/jVVFj7Us+tMNszHOCQ9SyyBJraChm5n4
peRCqIrq8/qN8irPfhlI5a+O9cTeh5JMpL3IqtMIN16KKTs6q5HZ5i1kkfmUSLRCyKsu14XRxf6T
lsHCl93+FGEwjbPIEx0mMBhl/mynWkMnn7A30dICWtNeO/S3iYrhsV+IGYVB0DlSpBUunakYvfew
YpoD1fCqZvGdW7yyv0rv+DcE24sYqwJj4bMG25TVUeaT9R0c92siqx4Y2wdWmMMh9UPtnqNvlN4F
nCslRlQorslyTdVKPHAZ4Pj6J4+fa5+cX+mpTDAoYgPkfYx7am5OGPumA58rFmPXPNtQQ5P5nfyP
GN/D0eyah3FdscdVUrjpWkQtBON1fHQgTYnYZ0NQXsMcijPvjpkGnJ8aaks8zu1o+vabg1pFsCxa
KJD7zE0sBOVp9wvpd9IUNdpOaQxrGU+YWWJ2AzXGuQHOlgVAztTRBwscvR7t8a0fXHgzwFubsNPE
SbAj4BrpuBUtC9bsb5s8QvUwORulVdFa0aWsUVEbFpxk/5kRRDMuv78dMde30Wj3vJ5nm4PO14eq
tjH0e1+7Dxq9gSamHgsbLQTsxgaZIGZj+w1bIdTGzL5hzc60qpHVRN2NHjaHye7gYrY4iSpMU7rG
AXquVoUPDfRkq8uz8/LU5cUgCs3m6Q30FboUjlXPg0Dgmxt3yOGcvJXpPFgbcLOjMebCdfD99sXL
lrXMxYDU16qdVfl2ijo9OZSgzWpB8l2nBDV1z7MsCH/E4SmWY43boNA59EeLjEZOxGhWy3XfwZbS
jUf09PSG5Jpk0cDYQzuEMJyMDvLtT125G7y2JGUJ4s8A6XCsuhQe0Lkz8Ccwg3WNwv7K30bqyj6X
HaBghZ3+FUvQkC382zjvVNjDWZDgJyFH5bI+s5CDg9AUQroxXCggAd3wsTv+kjPJ6ojNCyIJ51EI
xnC5S4liBLxD5u+NbGl9mRKNmxRyxmBAbH+O4GSkpczM2xa8AeB8eJ8rkKSC0KY7fMXU9dKL6PWQ
kOYA0apfdO7o8EKlxEzJjZv8DBGqQQpUZriDaRqezklZ302l1pw2OqEH+gswThmk5CpfNpEjYMt7
P42OVodOydBjv/W6i/ug50e2tzfMfMrWOvUhK8fbZtQMj4YuovSc0dQy7n6zuCpgXqcNYI9Avk4u
N/x7lFUHf7Ne4wk1AuFDskAMTM9Kwk2oDIx9yWEupIKywgbMeo3+VBpVrO3j1eYXCOexFR4coZZq
/YU1PQHCSt5JbiIOXG77+fanNgdGOWYfQOJSHttz+ZhxF2zB5I2slVBeJ7KAUZzviudQ8Ev+gXcL
P6bOwBx6KslLAS2CSAhH2peSb1BJT2rjzglcnrPxi05IB8IntkRSCry6HdH7N0fTv2A864cUNE34
7AvVfJX7bx9OdGm3wmHNHBKyEbTy3XFX1pO/eOhB1BKfLORxHv6oP1ZD4heuS+VIePMbN6Me4M63
WsWyw2Q2dfLXyJ0QZdTrAHDsaDWecQ9HexjeDVzXXwkJ3Ax9FnJM4NikSzujdzKqM7/dNdn++Mpp
69u02zMwLx3U75J3rUp2ROCA/wZCglaj7OlrJljQ7kvqIlJRTa0TibHLtB4JUXcyO3UPC2r+HJgj
ds2H3MK7wHFcaZ9UQNrDlUKnutPX8bHeCOMwHH7MvCoq5hacRPdnQfU9FDURhIvndmpeFVX/PAE/
zAj95XCqIrXlowmshkj16nKP6/I6ruC/us59noy6d63Rda163tRRtWypZyXvJhFZdIviH2nxrHdQ
mQquVe6DSgvuMuT1r1Q/Rh1L9HBJhBrBEcKWNOzgBnxTEruyyrO36oNRAPck2EVos0EihFsdb/vZ
BrcN4xoa/IrB3Uy31KwNmKvd2yiEWGwVV2DI1teJ5IYicIFspu9II3TUtbH2/kelJ43iZL3cAx0G
AuHYG/zILQT1f7EAlb28gNefvBgDk+/FcVRl9G8Vm+N904bUAyqmNsmLnfWIyRnzIiVTq9M/EUu+
S9HLeY3onDox1bV8ul1lm2tUuGLLpKNlNjJ+AzA0mDPjsyvFsv3OaOPUOOsRj3bC7R66SJI/3/JN
jZTDVYV5hmQrj+pGo18J+B/+KzP37T7q0SkRkEfHrjQcmGeueBfYxSOrPXkA2aZRdXPaE+vDWB4h
qXV9hOwXUoeHPEaJWwFXQG1FxlkqAzxoWJqQCrfB81EEyalNG1IavsCBBfCWYxNh4flYD4NtgPzB
zj05496W9NX2AigIGUpPZyIaCXsVk2OX9JGxuiuhZ4cZvtMA38Ekm54BnhUik4xmdUmO486umZUY
25WWzERm9nCCvyMfi6xhBof1R3F3FlTI08EpZxYrSVJzDFPbi0Mk9JQQalHtTVudS1iIaHAQChig
EnS8kAf9jUzrIGR1TBUsnbNsJrwt/rbTAVLAb9rV0Om9LVFN45R45KnLSOSDLHlLEyQIM+uRUpZs
UF+8fN0joAPxAugLAfVyL7lRrEats4QFzJ0KX6T8FRffH11zb5g2w8n8HQ==
`protect end_protected
