��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��,�y�}�ǰ�=4d�H���`I"��W�`r���T:tB�T4D�m�)�	1��I�t��
��8(�8t>s)ו�."[�漆���]�~�]��;�O(1#5�-� 偙O��QZ��~rL'�x[�i,mׇp���O�I43��4d�,�H�����SN��d���3���r��m���̨T�I;uj2Y� Er�*p�Q$Gm���p�V�`�2^���,hz�<p��l�Bxt�5��s��\yq���#�@W���f:m��T�	,*�񞭋����_��㧋l�	�\�:��uGd��PǷ��N�I��_����Tuv� ���us�(H�~�{2H�:Zor�Q	#%�3ˠ!��iS��95�,?�.���/�F�i{#���Tp5����Ҥ0{%���2vpn���X�����@l����3dc�ק�3	�Ed&3�ZN O���z��s�yxӡt��v*}ԫy nj#��lc��m戭k[��5)�A#�����8�!�]�Z�s�M���t��w�!��'ÒE�rv��Ϝ�c@<U��\tq+��&|�&X1)C�����r�A~��B�&�����s�:n{p��͠R�X⺂L^��R����c���f��J^?��ܣR�O 1�rV���:��T�4���AD����˩�F�w��)Dm�O�b,�a���1$��c��7t[i2>�ޔ0,S���󧇳Ϟ�ᒨ�-��}�!6��Jyv�醊�^_�(�H�(y^����o#����X��3-�k\8�M�T�"`R�DF6ȕ� �,5�;Ҭ C�k���1\������k�t־9�}���� ���QHF��"��t�9 ?��{E_�7��!����](�S��0�q��w�9��=�i]�1�GʦȪc�W�XC�|�$��}q�6����zf(����լml�dz������*�eLD�*�,�m�]ہ6����D�Gw� �g��' A��9�-nޢ�����`���&����BC6� ��\"/��D�,=�#��f�:���� ȍU���W0�!u����T�|.��@�}Id��r�����,�p���w?��� ���+���p�Ό�y]Y��tT��4���|�����2Á�9��{7�Td𚎕�l���օ��[���.���:�v�y����2�Ś�=	%�a�q���"����G�����D��y�qYMudH7ov\�^�
_��}T-Z$9��@�Hm?�)�rp�Kv�r��8ԑ�e���b#��X���<y�'��`��ּ;�m��:(_����w�-�� �M��<]"���>�i�L(�w!�>����S�#�5&Xc�~��`�E#E�����,y?��c#�ڻR
���e[8�w/��^�����������=x_��[o�Z��Ye ����}��'E >%5���XA?�+ �2+x��.�3�T	����A�jm_��x����u��E�]�=0 q4�\�ԋ�l��xsU��r�M�ި-�֒���v��ŪC�����Mvvq>d�ˋ��Ő�B������)d>���wӊ0C`�ñ��S�] _u�j��L)�%�3�Q��wEƳ��]��4,�_�8����Y�*@�;��1K��e����k_�B���.�4���WC��`c����{�+��{X\�"w����{Lˍ��k�N���`Y�JU�|]4�I��AH<[�������h�A7�g̼0J��ݐ!��Ƶ�P���R6�j:� ���vK�
[��E���R�3
��K٭���	l�g�EM����n�<�
��D>��=T�T�WR�o�/�,�`Sq�.1�Z�E�����la?�S�ڵ��1�X���A��/\q�X=�W2���/J�܃"O�n�Ӗ��Q[�е䅭Sy:��ϟHH�gK���W�Y��A�����(`�z
Ӿ���\�)^�]"��T��OҀL���o�o8�	[��J���iJE�t���M�4��K��!j�ߐ�x8*&�e��y2��ZyK�P��C�����'�H�C�!�=6;�@���_%�GR�ٹʕ@˕�/â=�l�?��G�'y_4FK�;5��5a����A3ɑã��JK��vWL�V�^<��Ew�r�r��õO�L�$!�����z��pΌZr��2"�_~���V�,�|�
��ٚ��?HQ���Ű�4>��f{�,Ti!8dV3C��{g�{d"�.�`��������mCo����p�k,��x�luM�����y�G/�&%�BH�1Ά��"&(�������I �~�qHpL�cR#3N��"��#�Ô�Qe�4@T�̅���*�xT��7������2����@�Q@#k
A���,�>����:�-�9��!z?
RJ?|1)�F%W/��������d��u��/֟t��R��5bi<4��z�Ђ+��B�w���>��C#�ྯAl���.?L[��.�r��[��!|�U�ȷ�mz��nQu�2D���]J~G�Y�+�w��;����
]�O��m>�9!�f�>s����z�x��]�wSq#�~E�ϐM��B݅�M��z��y�����G��Fm"��.��D�gKJ�͹7�|���VI��o%Q��Ԃ����+#nߤ�揤K���6��X�4���:y`HlH�ײ6zI�}�H���%PůEdm�y܍\�7��(}EE5.>7�^��f}�49f��c����VIF��<���
�82���0B�L>9s�d�ڙ�����'���
锁5G�AYu �*cdb��o���V���F���8ox�=�׹��t��`�sqM~����6��?,mC�� 8tT!�3����)E�clbd=�V1�_�6���	qJ��
�3c,���s�p��=�wul��̲�xW�8�4�8=��ϥ�\x� -�W8'�\���� �av����J0�)�)�1�U�$?,`͘9r�o�
�] ��u���+}5�ZtZ7`"a_�L�1��:Kc#C�Y[e��삞~*�W�����;<@t*�U`�PlT0<�4�p3�5�T,�*�V����.Ӭ��r�����SqY��2�����Y�ˏ�XQ������ `
8����z�y��8!�><8L����~3
a�RiǼEJ��KاJW0/@� �-���2;�؞7du��=���������TL?^�E[ً�1�8��Tp�.�������_�)�B@9=�e����@�-?8D���W�5�w9���)�	W?����{G�Yf��yZ�!ԩa��Q����`�I�����&M�¶姥��)*O!«k	\�P�y�c�ͩb5�
b.K�Ȓ��rq��$���)o���u��GdzV@<���$�ǲ����!<�绞Ұ6(^�ɍ��D,�g&���R�/2���^J��|�R�c�3� � *;h���TY��3��-}�0�4.Q�8�7	2m+�#���T��}�AZB3�"-sz ��|��"��+c�;Tj������Tn!Fq�_ƚ2V=%cu`��=�&�����H�Z�����ط��F���]�s��^:Zb��XG�N�ϲ!����h���䒲�JB��q;���y� l��-��j/�8��ص��"	�����Q]	��������<��-N�a�AC%3��B�d�����+��v��IE�������;N�IJ����9���9��H1;��^�Mh��]���� �e$��"˧��.65&����fjyM�7kȳ��[�6�;ފ5����8F�_\~���������.:�d�ҡw���X!5!��s��-�=�ol?i9�e�2"wH�qFr$_���lO{B�݆�.�`���I���VB	X$���Wk<8��^�c����,��o,:!����7p�=f�_���]�V�����M��S� �ߖh"��K>�F-�$����͹�>ӎC�Icѷv�T+���x56�(��i��4�/)�km�Z7��-Ņ�r\<7�uiW]/��3Q�wO��[��CM�����k�c/��L��<�L���2�	Ñ��{�4*��f�_$�� ��B9v��Y�����M*�o��c�����IZo�2h���Z��}�S�C��i��l�X��x�ju��6������n�s
n��b���#��e�ߴfO���0ʠq������f+�&�X�!�6K��j�5k�*�:"Hʁ;R�	vU�%�(�;��-�x�k$ӄ��#A���k��F��w��`��}�I�^\ެ/{��u��򨘵��DɨV��$������V��+mJ������"�Љ��[�Aq&�$�ܢ����6���V~|�j��fGǹi>{��/,�t���Kk�r�gꟄ�J���9j=�Z��,XﱹHvʬ}�	w"7�5�U�;X��<���
�V�_fъ��-ׂZo@���oǒ�.c;Gc���5�f�v/'� ��5m��Ҭ�QQ���V�w7�c"�[p@F ��:U��z�k�h��@y/�<�3y���������&�j:�z|\u�<�{�����$*�z��+|�r~��KT�	�l7Ъ�)�T��y��wb+)N���r��k�8z��?�g��dg?��1�Ì���CV�C��D׶��g:�T��Hr�yX��6Y3V`�2m�\<�e � ct���w{,�
-�
Wb�i(1,W(u��v��7����|�^�>�1ҸZ��I�ӯkQ�⇯�G�K[�a�ů}��u��ܘL�eJU�%ϱ4���ʴ#��|��!ʒQ�d�\s���N��D�s���1�þYP[�k9�h��REc�k d����|�Tm�ΥTZC�s\�L��r2g#ɒ�ɠsp���;��<��Z�Cg& ���_�4�G���|�E�[�!	5����뛯fG ��A_�5�PU��`nB��Uz�}R,Ik�j�e�n��|�V\�d?ˏ`ۿ������4��^񈽻���h��Z���[��m�gw��0�N5A!����VQ4š�U*Ya3��y2�u�/����0h�;n���Gj�q�<���ч�|,���&l44���R�H.������E;�̃� �:�wuzZ�B���z��v���`���JV�['xEX���vF^�1�ܱ�k�a�uE��IsL"�ix�y.A�@�9��0f6�/��1ÀCK@n�ZJ�6���R�N�t/{w�!x.�SO�Bq�sro�p�b� ��T`�pdk���S���x*�늭�W7B�N��v�huSV ��8n6
d�C��@�Lt�7<�e��`�jK4�N��o�*�ǐz�IeH�!3�5I���͉i��n�z��o�$�ܸ���X�t���$�b$��2�6���3l�Y��W"o���ef���o9|^����:��V4d[T1h*8�o�/8x6[Vh�a&%|L�|��!�[ߕ�S� ��.A���X���@rǌ��4"ّ�x�u�p�V�$��C0A��ɻ<��ܐ>�N�-
�R�	��0�50��?�����ʳ"y=�R��$�͇e���1����*7PJ���wz���	O�Yg��a��8dg�Hݤ*��}5��yRD��ߤ�=��+�K`�Th�D��D!�^#��*��p%l����}S��u��
��� ��zc�QP
��lsż��q��XQ/��2Y��0e1����/��9�D� u���yJl/]�*w�����Ħ�7����'mXS�8�dD�NI��}:��р�c�)U���y����*&V��Pk!d����]��_y|GF��2}�,(�ؤ�g��&��}����sJ�sm*�쮛��DS��P5���wD�h�j�з�� �r2��k�G��M�;P��և4g�=�k�g諄?9�%Dл��2?�K�c��M���\97O�2��9�µ?_w9^��*I��Éݲ�*��=���A� ��ʦ�����x��]=��Q(?T&f�X���kx���H^��O�Y�LmY\�\�@�A�f��������|(~��B:qZD��<�7��T/��9l@w&T�`9j��K�Bh.���vx���R���z�˓��8�E��Рξ�Alk#?��p����'����=]��G~hоv~��o��c=?C������]F0T��v�E#�0��;߲���3e����ȩ?L��f)��V�sD�YI��Av��=�Gô�'�H|7W|���X�#�KKm˦J���!��\�[�A��������r(�2��Aü�q�g��Qwʝ��r�-#��f}�_�%C�A����O���(�4>���R��u�@ُ�c�^K�0�����%/�ցV%�F��u޴�2t��m�DV��E[����D�M�I0Vk\(эB��K���K������@3�D���_������ �+��x���9�Zf,@4խw��S��;��-����&�`I�/<����g��k���%u\Ni�U����Ja�m�G�g$�d[^ޟ\������"A�'ar�3�D�W�`�Kr	��8o�L=$���n�\�H��N��9a������J�9B_�Qk��az����]t������>�`�C��#4e���@7�؜�d�	��4�[�t\��������?z�����5��>C`^�����P���#�T�E�G��Ab�;�<d"��e�C��pgm7mx�R��)%G�C���;�}_��Ar-(]�v5�*�{х��i����4L���~��O�wQ��#&���Z�I
/����S3`K��$3��^|C3ZP��mK�Q�W)��2ʫsz�0��z]xTXE/��V���3��,s�&�q<��qV�Aj#�d��6�G��Y54�|��L4Z}�-�R<��#@��F�t�:�d�-�q�o�,H��$\z� g�?������f*@��W�J�<������Eq�m�@�[��Z�= $nicu������&���5��Ф+�\eE�������c�1pI2�^=��4�>S�Z�������M�Jt�"�Ej����U������l����Ս%�89��$%�[:�̟��řP�ꏞ,|$�[;�N5�����LF*��Ր��d���;��%9�4ak�1~B�Xh�҆��<.�j7+H������R1�L8:�a���C�W�P4��˿t�k1�}0:�ل��N���&:�yq��[��͎�|]E�ocr�T���n~l?bOg��/�&������C�;dă|����Ba�ޞ�M��gk�]��(�`@�p�Q�D��wQ����@-='��3M7���Xb�� �����p_����]3̨7������D1���l���Dr��RsQLY9���+�:N���� >U#���?Q��'��H/	�(���*d��]a:�I��d�'�v��ƫ^�y�������(P f˞'�*���݈���o�y���,=�A&}��n����A�c�_"^6���+x��?���*������4	
H[��^ݧJ���Oc���~O��;*c-yoT��Y6��a΀�RRsz�Õao� ��PQ�x�����TP��9���0+l]��?�j�������+�����8���X�㤠o߂B��Ae�q�Ͱp>�&�d�z��������]�����)�| ���w+A�����]�E����Xk��nA]��4X�b���.w�4����j���D��?�qZ��5�#�#6'�j�\�3��h^��V;"@��A�K����i�p����9�7��c#�<�-�N��;ˎ;�5L�����z���#��?����;\f�M�8d�F{n�O�[��n��Pb�p9S7]bc���*S��h8$$<B6� ��p٘}YZ��Ҿ9E�����b�Y�[��
@��m%���c�ku8m�y0=���*�qo����>���_A��@Cq�HL�[�t	����
[��|䦞�����D�~���<zB?v�Yݢ2�x������8�m;~ ��l��L3�*=��pg�"���&�)���E,ظ��<��Ď�\qۺ��um$�P�"���&_�O]�R@{Ş�:X���ч�M���(OU*�cz����"�Ra8ϟ%?������L+�b�$6�:>����#�Z����?9�w����n�כp�#���v�V�JI���bP��������M��ů`觞o~*;��;7�t�8 }�Y�a�c�5�%+�'Q�plu�,�]L���M�\���I=�ܴ}&�_Ya�0�xz`ZF�W'|�l7G����ܹ�Y���^��洑9Z�h�P�V�K�0�Ԑc���~L��s�0�m9ҷ�>}��6H��)\�Oc ~���k,eF��:�8�J�P�b�`D�r4K��ͦ��:8���n���G7�a�D��qɸ&��iN�Y�=$��D�,z�C��_X���hS��#i�D�$�i���8&{7gL^������42�/*�n�9+��2�$���7�ܜS��G^�7�I��@����9��EKP7�����a�����zN�֟fx5)w8��q����i����P��G�I7�Nyv�^����n����T"�83�'��@�~������m���i+�5`�`;ܯ������l�$�n>��7� ]u��v'hȪ���<Ŵ���Y�&�����?�EaD�ż���܏���iO<�d�K�,d�Zk�}��'s�a�,Dn�8!k���4����%���V7��4�5��m��!�m2%;�I�A���S��T;HX�T�*��2Ź('NTU�`nƭ.:�>F�?X�F@��,���n"��[sx�7R���j ��@�r�
���?������-�ٞpE�@�T�jE�	�;�cw�b����st�����Cc\�%{�d��1��n]�0�jI���[<���P\�!D�����+n��ѯ'��������<��y���=�5�6y��I���n�<�����B�|�;�n�.�i���y� k���.iD����ЀE��[�m��m�?�>MG�\I.����}EY|\%����5w	�F+�Ž`rǌ�$��,Tj����bO�2a���|����-I��ʴ��d���r1V���^f�N̴��ƕ�OsВ��$��:l .h�g�t�˖���۾C5<nbUZ\n��[$�c�������[���c��W[�{�+�%�m���K��ǭM�F]�.��UK��݊�c���k�N�2�eK�����������H��BBM8~�E+�f��$'޻ABf�yS�E3�qY]�6��Q��6Z��*�U���;���h�lYX_NB��d�I��{-�����Ғ�40��49��M��̻��DA�(W�����$�:3!�53�*��HT]T������"u396�I�߰{��ի�*q�Hք~͗�3iH�l���at����9��q=��T _V��m-��zq~�/(r��9㏯\#[��q�6 �G9g-�>��Ĩ�ř�A���h!'Sa[o�L{*�_4����[Ʊ��b@�HoP�S(�c���Ķ=O�~�!���St�/��U�+�磶W6�k�X0�V+D8DM�j�k���T�O1��ZC�j�-�C�Ĉ0��v�\.�����v� ��J���Cs�� nTQ���-t�yD�ljY��Ks�+�3oz��0KI�<��;���G��m sO�Usc���:��8$�y��0�"!��K��%b'�m(�D�Q��iYz2�&N�F�N��ƈ1�Қ͊�I\v<㗆��5���??Y�;h��ǣPy����=+�V��Ѳ �A��5dx���í�}�s����z��p��}I{փ+ϤM�9 ٛ ��+,�A��h@:���5ظ�y ��ltP�#�6��&�N�g����kPP%�J���
lf�����Y�ʤ�\�H�R{|��k.���+��e�������O[�Ŀ=�S7)�hg�c�ў�Ѯ@�I���G%߷�]]�u��^��;�љ�?���JM>�E�Gv&7S+}E�������Uu� ��50�_r��Ͻp���D�dSs%�m_�@C����	بAݍX_Z����Iy6avEA�P��zf��6!���R����ܿ��f6���-km"��H mS�'�x���4i��������a�#�I�#�QnB+�щ[p��7� \�"%㧂�f8�d�,� g?���ٳ�U��aD�����T4�F��:�R\ґ8�$+�"Y*�_�.]Q��*��t��w+�,u)�x�U�W�h(��e<r��b�����+ˇ2�;�/>�ͦ8%�|=��y-_�J��YJ���������[u81�&K��l�M�ݖ+o�EC��<d6�
����D:iÿؠ�FCH�w��P����ge��L:Ap3��OPU��d���~�=��T��ϐb[�������ae��9�O'_e�'��:ܬޒW�F�u���J3��?�<"�� ~j!�dQT��Q�/������BE�e��%�����,����h�J�'Q)9�l_�aá���8�'�ƾxF
���.�U��_�J=.�3Y��r�l7�ȣ��\�Vta��Cᐶ"�!/tҏ� �X��ͧo'k.�Nr������~�1N�ߢvX���Ȼ�?�� %�d ٴ|��M�be��Q�ܼ}�ս#L�)C���&��a�����$&�<D溮����G2�[C��yP�	\w@W�k-m�Dy��S���E�]��M�ҍ�R�s7B�1x��̬��l	��#�a�k��x5s!�[�ݨ�E��
�]�H��v��Etz��ѥӟPR��^���w��o�C��wz_�������?���g�a	�qC�u�n�ԕ>����ɋ�����ܚԕ�/���o��<�l̸�oyu�55ܶ,1)~���$�΃G��b�t=� S�C~��O~;w+���wY࣢�6ٲ�{I�F<#��o��;�  ��"�ٵn�h�#�R�#g��jA%R�����+˅�X�ǳ������d�vh�7$�Γ�Tذ3��U#�j�&� �O
��-W#�"�����Q��R���w!����*�L>~|���K��_�=Jl�9���-�|+ n�����t�OI�ψ��*Ŏ�X�^�����r7xPj�0�^�J�}�|"�4,�̧m%p6�gc��@�#т��3��Ђ͚�3<�\�iM�30��Lc�E���rɺ.�����𰠤�m���J�6�6M]�[8+-�j�St��Pg�Դ�X��!w�vP��@
-�������i�M��;�Qy�GPD�8nk"߿����"�$�櫌!bF��R���r�H���?�y}4��r�x��N�HJ��)�)�*��f��KQ����bq�����!#i��ýGТ�ru���h�}�@_��$���ޜbp�����8���:���䎆J��(�LI�� ))�K��i����D��>��"�VF(ҡr�+9=��5��v^%�-�|2�:h��1,�ݿ��u�Kץ�ە�g^�׀Ԫ:=ۆeG.>6�V@�SFC�1�l|��}� �����	��~�	�q�˿[�cO�$�L�I6�vD���s�e��R�o�&�������µ����.��7���f,��.��Kg+L�J�O	Qx!�1�IxO]2�e�>���^W���[ި�V�R�Fl�+�$c�OӷL�񁵙�'���|^E���{���R��i������à�bta�[]^ܱ ���K�tg4P�t2D_�s����eB7���QH��ae�����}Q�E�'��B_fb�C��o)���;����Z�$��_�'K��	0����%	��K�����_�v��QY�U"]Ѵ�7.o��)QW���Ǆ�7�,P�0�D�bwk���g����F��m�Γ��5_�����v-:���u��@�i��s����fzW����#���1lF&�|q���g��W��Dw1��H��l ��I��t))6�F�&s������$�
���gHb�����o�f�A]$�7���O������0�Ҧ<�~��;Z��ɀZ�Kc�VVC�b�� �6S�w��$$!w_�Mٱ�:�Π��EJa�i��hG}{ٖ�#�I��ecĂ�{"~���:aTƼ�;�)�ξZ"%/9H,�'$��㊫<~n��E�.����c1��JW��Έ@_��,D��=�E�){6Ź�҃[ � 5\pK�z��R��p0���j�BɆ<��cZݣF�(7	��k�qsc�ؤ�{�n�h%WC�����J_�r9n c���|���o��_	���7`��C���%u�h��F!R���H��P��_�gA{c��%��������^��vc���;�ޛ�@���q�My~ځ/n�����|��\a�Ho�	��(���l��a���(�zl��ȫ'���� zN����]�~�4���ɓ��K�QR���U����T���o�3�ܳ�@ ���W[�������+����H�*>Ѵ��Uyg�̍<�O��$慔B2:�N��{��B ֏	�!P��������Y��-��1����-�WZrr]�7��&��h�qvw�Y�3��>���ts��V3d*��C�ȣ�����Xœ�[�g{+i7����҇Z+�m�Z�
ܘ9���1�h���*w\}ZU��-� ����_oƱQ��h9d�k�����A�o�k��2c.�I�����
j��z�`��U�n\���u_�{�Uqo�9}�����S/	ƥ�\��Qӵ�A@�����8���s��-��>�%%��l׻��##a�jP�QF^i8������<�h�	iT	���,E�̸�t��A�r�q�\�}���A8����m�}�<���Ԡ�v,�L�����A��zP��e�I��f6��_�I�,|�X�w��[	އ�3;��C()�ڝ%'�n ɐ�m+���f�f��T�����RE}�2C�T��g���e����Bc�N��Pc��;h��3J���9��+�/@5P��ܐ�M�m=bl�%^��<n�<��PE�$%�h�E���� m0��v��v�d���:�|�@��Es|�l��L꣖`RKX��؂�����)ԋ����t�%x�.Ko�yxw��u��O�|8�K*�C����U���:Ե}p��]3$)B�ދ`��J8�������N���o����-g)�夭|>�2�z,��Q�wR�FxJč	�}y��^����5XE<������� x��� ��]+��M](�J\A����-Y�q���L,���Q�J�I]�c
�̶r!���'@9i[V�/��p/����臛c+�g�i�` ��x�u�X+e�P��DA����	n|�Ű|Y�t�5�w�Q�,��.�7�$H��Q���9�	@ĳ8l����?����ȢQ�{	`��X�?u��Ң)w]Y� �� �i�د֝&��2Bl�)���h��cX����ӭ���YM]lZ�uM3._M�"���2�iH,X�8/@Ip�e�Ո w9�c�"h���[�� 3�{�Q��'WJ�g�eeC�����%��G�Ids�v��&BvX�̆*t�/Y�'�XT�@�ۖL�QN�&��:����ֵ/�ٵ�"\���ǆKR�]�wA�k3Y��/�#1h�������.!����;��QQ��`�Q��iZF�{��x
�"4]~�a��؃��T�3l��s2���=�͸�DɒL�P���rE��'AT���+�*F5��4��Y�q%�F"����2�,�* ��c�ᓕ�yU=���H��W��U?�_�u�)JtQ2�!����I$o��0��܆�����=Z��(��f���l�V�&S1<8X�Y�0����;0���\�����*��{&��Y"��e�\��sJ1�����4X(�]��H�f��������b����A������r5�f=p�Ϩ~�W�}�uM?�%�U��н�T�2qs����#���LL���3�S�J�O����;�>;S#��XDW�������;U[cq�TU/��e��dswjP��+�]y�B��u��\H)�� ��f�i����,f{$e��?��` o�}���ݯ�R�gg4$0ȡ1ZgX��	G�9��������^]�Wkq��t���MJ��������^�{��I���e�yJ�F	�\�JE��Kl��!�݅� ��"	yc|���=����LU�s�����K���pr��4�b�?\��`54l�8��r�y�%�7�����  ����9q0�6�E*����l*,U��qX�D��