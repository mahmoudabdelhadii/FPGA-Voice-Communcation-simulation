��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���/�����Cc��<Nb��.�x{�>��0����=�����=8RLG�h+OLزV����ݗ�@��&�K��4cbXu�6@A��?��I�=��O�s=���
�S�i\��D���d3�q	��9/�I�w`W?ދ�S"K7��5�,l��C���
@E=D��!
����荾Z�V�h��c,Dt��&�����]4w9K_9O�=l�uE�w����[R�\�zÚ�-J�$����åCj�[�
����T=���K���h�����,������#�z~��?�G���B�~֨1)��k��yq�$/ju�YA9��SX�{@��mWt������w�F��r���������O)�mC�&�����$��^_��|�����=������A���_"�s���50��-�ݡ��kVE~�cu��'Ah%�����v2ݲK:|�g���7/��=Q�u�~��qC���
qSa�a�n�m(�]�h-�FK�]�Z<��K�b�s��'�����C$Yכֿ��h|�[@lXJ�*Qm?�аR��(�v�vlr�j)ڦ��0p�s�bv��jy�-����(��N�vהS��Y�n)!��\|9��;#�o:�#��9|TWL��L2=�'���$ƫ���19�?�:H�A���T秧���,rJ$�p}�a�ڡ�rn#9���~�1e�[e���!������{�T�7���O�z�������쉎�<o�j��D�7��lS�ƃ���F�V�:¦?�,�:4I~P�o6����2
�ԫ�#��G롔�qH���'> x������>I�nN1.�yφ�V�ǹW�)��	�3���k��c�Rw�buRA�8����\��L+p����rw3v�FF��8��Y��8p��s3jL&���9>��y�(r�I)ռ̋����̩����\Yޗ��L���o`i~ɦ�.¾���O��HN���N���#�(����wC��p�M����//��l����3����&�]?V̵F�XQ,��`�~�HTB�<�k�� #0���h�-���s�ӐXY�XO|������v��B��q,�>Ip��IZ"+}��}�A��I�L��,`+��k?%l�_��<������!`4o ��siYSר$V�=˘d��1A#W9zkv�aP��
���e �T����h����:k�Px�y썍8��	�kF���B*;�!����?��9�H�DNK���*�@K��Yo��&�.�NX�����R� ���}����Y��؆&t����"N[�r<��������5G#j��ᬡW�-��M�'�j�S�to�X���F���Y(H-��<�/^��Apk�F���>	�bC\�E�2*��6�/��;��8�w��1�����ٓ/�)�,R��\���qe����'�Y��s���>���S~E�˘���zG��ss(���K� Ad���ru���i�0z�����a��Z9�ew�8��>�٥��W(��Ɠ�e_�&���g�� ���~Bt4;���j�D�[6��� �^/=��X��^�����F��?��#�s�OR^���G���Ys#I���9F��%�q����*̘�o�W�!����8"�F.l�F�,���<�����SS�@r#�J������8���I!D���(�l���rI1�VO���;��r�4`�G'�n�J���HC��P-?��π��躘���?o��3��R]�g඘k���o��m�&35��N&�����$�AJN�����Cp���vĝ3]���/fI־i����3:�k�)�V�D����\Y	Q?i�9ST�3�=@6����*^J)����K!y�b���u�u�[7�E-Κ7Ͳ�բ/�*Ғ�Ӵ�ⲃ����s8�b�����9F���d^t-�Opv�]L>��Q)��bӽ��e�,�;�Ƌ�'��Q֎�UT3�Q8Ӕ�ʿC����[\�J�}^��M��KJ�P��b	t5�tMv�_�=���	�8��R���v��>/
Q1��w��s���*��'�R�}^�8��E^�� iE�>.����YXN�ʓ��8� KL�#��;x�g��5��:�P�X��EB��'^t���B^��ӷ�]�-�&>�_�������;�<5=>���W�3�U�9;4�g�j�л-���1�)`��#�5�c$�7\q*��vksd|�� T3N��ob��\FU4"V:R.v��5�騜Ix�{J�?$[^nH�ڙ4J�r!�u7���+p��3�=/^	��Z����(,�J��.�����Ë����^W�^����Sh�N���Fc��C���t����h�W���Zc��%�<%e3������$���g��O�w�FY�������١y;�I�%��u�{ JNnwյx߸��e�1`m� �=��h��z�,�6�YM���
�'�b��#���L�R.���~x+�hF+��]�:gG��Cx	s�_��/J�0k��"^�0W�� E�^� ��έ�>y��7�ų��t�Ѥ��kL�,:1��>��u6kz��R�g�V_�Pq-]�W�:?m"�-e������Q�x�镁�����g����^w���a��_�2| w|2d4��;'*лeH��\.Y]�"�*��λGTڸ�ݢwGhx[7�'��܄"�M>R��V�#�z��M&�	
6�*����(f D^]��	I�|kׄ�3��:�y
�'���R�.���~�����"��FAP� ��zA���2�m�3��B6�~us�퉃�]z���	�?�����)y)x�^ )�:l�)� �}��S��'ş�b,�a6�s�����bh%��^�po}�_1���ϑ��w�|u�H��ϩ~���!��lPRZ�?���f�l߂Ho���p�ۑa!��c�X�q��i��kf;F�B�f�KYwitKg��w�Sj�x>�� ���@�Z��]����r�+�����y�LF9�%��buX4ot�5��ڟ��|zʟ�bo�h�M�}���%BR{�tbT�r�R	�u���Ň.��;)�7g��O�żN�d|M��A��\���²��1R�m]W�Њ�����x�edm��P`��B����6�Uڦ����THO���\~�&�{��`ԏ���p�rL�<±�Nv}��=����x(<֙ ;�|Ƿ�Ai<�M�wˌ��ƬdKs	�֔�V�Sg��Zs��Rϕ��0���c�$�jm�_����H-^�+��������.lʬvT�_֬
���Ғ���?�5�p,�΄��?L;g��n#Ǉc�}�o��C����4�{ѵJM�i�`.2tܫF���\s�`"�Ʀ<�8��+g�wq`�W�J���`���.�Ӥ�����I ^�`�s��乌PK[�pr�c);�bP�c����y��M��}�����ڕ��j޷h0U��4xbB�>٧Q}^����,�ת"�sS?aԓ#2�B#g$�ZCa��\��!s���j]8t=�׸*��i29)Qy䐢��_�Y��Уa=���3�ƅ�6ˣ�}����-����Fޙ�s��!x�)��&4pBpx��/fB���#�o��+Z���u�s)n����Z�S�{�9���kaWE���5^j`(�Q�G�bXT|�ωU歵r����x�����r�E�*8���̈��%��$u�NUd-�q��5�yi`R�eQW�'A�&$BUu[��0v^���;w�3=�o<$%�cY8Y9�)ډ�@���Q�Q��2Y��̨ ���J0\����+�= a>4�!��K̉'��lMe��&�T~�">\�=.$������_�}r����Xe?�z��՗C����N1��KD}R+�Y����*���
A0( �{Y��@�j��Z�(�@ەD]���>]x^����~�זk���G��6���]��w��5�_k��f��Juό��鶃���
NK��z�υ���B�1�lP/���eņ㲥�	-���wѪ��=4��u57~[V����<9-�S#�y� oޡc�;<��zyW���,Xr�t��pk�rp(�q�_r5T��J�=8Z��C�e{π��_5tH�jGi�[��}ɣ��R���H1����LE���g
�~���3%�>�Bz3�A�ַd���a�9F;��d��j��v� �6���`*����Zމ��L�"�qǻ��c�ڗE/�����@��9���wi$w�<�6W�t���C���/�)>�nfgT�ɉ'ѢQ�T-����b���C_�����C��'����³x���+PC��ݍS���@����S����GI��i���7ࣖ������f�'�4�I����c���J�SڃlW<�B���&����*�#��ސ��|fD�=FW�$����n(om�P0���1��`Qk�s����!��ʥ|���9]C���Ǹÿ�g�CI]l���>cl�v��m��rU�!��@�<(�fC�ot� <k��LL6J���4�'���Q��	 g�o�lJ;�9	�OC�����]��MR�j/�\H2G�� }�����l.fJ�'�[e��2b����I0��:{.?��Ǎ�w'��Jr�B�aM`��O�|���"����Gj�)�^N/������D��l7`̀_�~�I=U�w�~��F��u�n���D3L�x{P[���>�l?���2��ҤZ�9��D&�"z2)�ٞ�5JtS+�KyA�x`b�k��Hl����ᩊ��L N� ޷��LrNަϼ[<���2����[����������N��R � %ۼDU*�m<�ß�v�`:�^�}%pM��C(�tip�3˥��
nDe��ر)$���b�V��&�o�?X�eI�����^6����x �Q�9��n������He>��4��hQl��H��!aA�`��FIU�#P�k��.][L��d帪ж/�@�ոC -��k
���6��²��3���P`wH�l�0��%��JK;�v89�9_,
3xi�q�D�	��i]�5]v%�<'���(d�{jb����2��!(��I�"Iv�V�s ժ�jψ�!9F׻��:�!�&R�R��,SΑ���xֻ�jP2��_��S��wQ�KדwMłG�D���I�mv�x���̲�M��kq.(��^����=���ZX�5�o�$u���"�-�)b���b�/�Fy+Q�1O^���7�НL�^J�\���mq9�bZ�?i��#]M�s3���vw�
�z�D`p��	���۲2['U��!�'�7����Ң��ױ�%){�$�[�<3-��}���@�����l���@�=+X��/�X �����ȫn�	���<d�&��0i���!�<�E/;R�a(.��|�Bg0n�����	��n�ވ�q��Ie�s׾J�c� ��NK-�$��Y[R>P���%���o���[�4=�J��Z��$�2��ϋ��J��?�m%�
ܞ�I0H�{Зڝ��ױS���RӢJn�ҵ�g�nO�b7�����y�ui���MҪ�@4w)���GV���Rc��)��4#s�52�mt�*I(d��U!Ƒ��7s`b�����c�_�(��|Y�;P�_��J4����-U�z� �y�0�'S������Mݗ.�a尓�s໯N보W</]$dm�͛{���6=���(�Vy���WM����u:Lu1+<d�-.��S�>�!٭��T;��ӿ�D��z��A�����*۹�4�d�=R!싔:qeQf�RLn;}TApmB��2x������� �B��I;]w�b��U+=h+H��Б�گ�H����!�B;]��<<
����d'�����X�� Q��2�>(���,mi�~�C.ή��/LiZcK��4��Xu�P�V���b�S�B��=����W�$=�|u�U�形2���+J�RE�[-i�}��ǈ��x�DG�}b^`�'һ�,s��h]�lH�=�W�AkjPS��\T��h�*�/���#ذ>M&
��MW��&v�!)��W����o���{cTS��9��.��#�"-:D�8�T��2y��-s��S��B��t;��n�Xz���̼9��J�I�_%ځ�-��d�@��� �u�[������w#�1̞�FzdL�2���\�}�W��YZ����+��+�5� �}`�#K����N����������&"`6�kh6M�݊`�\���h�-~J��#�/T���׽���{WA�Ԧ�|���Ř�E(f�� ՀVl[2���86a������!)W�U��c����
9)�h"�ȝ�v{���h|�N�k��B߾��x9t�̌R{��|�J��x�����0���>��S��~Ht�D��nd$s��Vt�i0�F���ޠ|�xl�����VM�����H�E�5(�P�yQ��2��"�7?�B��M;���;soR��,��X���e���rS��pP׉�\��h��
v�4�$��֘���Ή�p���_Q�\����z;���.��{.~�1��Mq,7�0G{d�Zl$2����Wz7��Ɯ�[���˫t��Z�F�j6��W���R_���N�s���qY����'3+Œc�1�'TΔ�mG����(*�������|���{8HJ��Ǚ9T˯��9�I.�
��84��^f=H�����N�d�s91�ڛ�U��N+���ю���/�J�.M&��
�.��.@�]�0�E/r�@�<ᖐ�9�N��:j]hQ٫��]/?�x4M��`UD~��M��F�����m�v�R�[4O��$v=��:`�]����k6�D�~`���%����{�{�
Ac�]���`R��6qE�!V��#�2򍓒��Ɛ�0�~�3�J�y�0���.Zv�$�1���;��L�������}������D�>�z@�:�=�ʉ�tp��Jc��Zpkc�������
�>TK��k�kk��P�j�6�k��Σ�o̦Kf84o���?e����t�#>h��[d�[�1Ӫ���E��x����%�SG3�~���
3Ұ���%�Jם���z�^��?�oN�&��P����d�ȣ��,��7��.���q���d����n�C�E�2�����h�Yҋ�	����Z�I�)	�*^=���ty(����!�q'��RV���Q��B�j�L���~�7T�/?�L���?4�)�Wc��8{K4����q1��u���F�����Ddˀ��oz�T/G����a�U�)E>7�*4^��s@A�
�T�m�ϡ}#��i�GaI��hԷv��e���GA�Z�IG]��]+.�X�	y4����z�����{�{M��3٬)�=U�A-.��+�m|��wImD�Ox�6���g���O���DO�W���z٤9_Y�H��X4�	�d�b
�{�P���`��BS�׽a�Zh	�呞�j
sPO]J�\��Ѽ����q�8e�Ȁ<5��ק�� ���^~�5qss\���Y����3�e����*|a ��ߖȿ�!9��<���3��@�ұ�{�H���!��9��?���b;�p�4�q6���sܓ6�ۖ�������iG#	�����&ɨ,Hg e+��.���W�O��v0�&1�7PC���97��� ��C�q�ҭ�����B���I��C��+λ��y�����VO����!��~�����)��!l~W�O[�-c����	iYv6���UVÙ��4����t�[%��ju.��^�'O'�>$̑`��OJ�V@�5��8Y��T�EO�!��SS��lX	�䠬�;�tl��Q�)�q:V��*QG���)���Sȅi�_�k~j��o���3QC�F���U&&$�n��d��# �|}�1=����Ek�t���0ф�xamڂr�X���\ki�N��D����Lș�Z���Z�o�D���@��#�+{���u�)��M�d_��is��{��&X=�cRظ(G�,N�H���G�|��A�|������	��La�Ť�
��" �H;���\J߂Y�����IA5��[��KM@?ֵ�ea���6�S>?QE��Ͼ�9f�v��Yԛ�oM�}Y0��[]���\���S��5��c\�|/��,}�Y�(���})����\��펣���4E�D�ل�lm���W����n�y�=J����r�`TN�ќ/���12gF֐���� ����j�qTM<��@-+�J:]�^�U�*���-�����%����)<6�~ W��26�_�ؿ��,DQ��bXqX��_�@oK
�ʌX*)#<Wa���9�Z���^W����29�)����6�M�����$���lG�	{����C?��<\�F�>�V|�f��~�E��4V�	��9���"��E*��ܱ�] �6��j붷��}���K�ˈ��:�'hf��Q��8;r�	�(aX�s�ԽݜE�͕�pR������z@�.;v�ɘ1K�{]�����:�kl)�ͽ��w�\Er�p:LW�Is�h���z<f;l;�R���Y�tQG~P�@��˕����R̿�s4XK1!�����'�����S��o�[e{���`B'���ֳ��W}IY2`,�ݤ�@;Q0��� h^���<�I�h�����ʏ�Im%��*(*��e~hH�uKP��#00΄�^K�`�Xve)���������X←�e�\X�,a�f^���c)j�q��Y���4J����A��v}��(��+�Tλ�Q�m0�pj�f�/C�ɪ*m4N�(���u6V||��f�Z!�>�L*�*�4N`����&ý�u4�U��<س�g!`!]���:���ê� ]�6��Jǜ+�?Q?-s/*�l	����'X'���1��5t����~��NNârpL�/a�P�C�f�����:iRh��%o���ȋxĄ�~rX��L�]l��]a�^�xͱT��cjY�+գt�}9ݬ+���Ϛ0OZ��E&�7i���_ sj� �\���@����\[R�̀���L{;(D�S�U\�vcD�V����`h�����p[�@��ҭ�
�������_��x�F�}Xe
�����_yP�4��rD��������Y�c��N�<-X�:��3{���F����/�6ÿ���1���%o@?9�[�z�X'�D�|s��y�I7�$B���i��������5���l�I-���t�Ye���ZR��vY�E���8[�$�K�)�����᩠M%Ju��S���_���2,l�����@�P<�zS��ȞS]K6̔卞XNʠS���e�d_�Hfۍv����13+�6ٝ��Hr_G�㔶H�w��G�}��Ax�5����N+)���p��ߡ-� ~���r>�O�[?5g��A��\^�bz�d�+<�?[�i���*���p�ydH��6�Z���-����v~�?���}ۺbfQO�+�|iԼ���j/(Ԑ�����xm��������b�7ȵZ����2ұo���c�H�ށa^ K�'��T���#D/s���,ګ���9�þ�ϕaCQ������n)�P3P��)	U��,M�*d'N�(ϗ�����(�d·�c�w�J��V�;��ă	Oow_$#��S�j-��F{��g�TdǢ�֙��q�٭����rI�S_|����-*}2��3z(bi7���6�"{��L���,bM����#�]C��˖+�~nӗ��ѡ
ۿ߀@7��V�m,���a����J0[,��d���>E�-i�����ﮝ�R��B��vv\���b-�ߪ�1���C����0�G��94�4ݳ���s�P�Q��v���K}#?R3�� �����1�K���8w�w���m��u8�1�{��S�Z�5Hf�R��T����u=e�| �Vh���u|����9때K(����0�@�#��R��,@K�;N��'uQ��A��������������[N����� ����#0`��g�	�ʕ�<Ÿټ���DbH�'B�Ԭf�����9T��X�ր�f�EX�Wlф���
�%�����V)���O�{;�����?���a�v�o��-e����/j�|*Q|xlid�aJ�18l傍�}^��;ȏ >W<ф���eIl��%���!c�E1�iyك4���:ѯ��-T�j3EK�>��_	 ��M��t�4N���t� % u6#; ���&)�ӫ��lBR���7H�٠�{��~�$�C��@��Ε�En�؉֧�;�Qޒ4;�~���aE�v� �%ɳ��.�Z�_�40e=c���;��ZD3W��5��Π�%������6%���>�-/�O,z���oЊ�{���S�l���u�x�v����sŷ��U�V+C�үH���=i�>�v�J�ۏ��,lL�ͨ�^ۖ�ͺh��!_�$�f�ږ�R/��hwZ0�/�J�_��rV=��+���*���+�Ik�!R�
�|<Ey���ڼ�g僐�c��!rm�;�ܒLh'ԍC^�m��.�Ex[��H��P����"��]�����+ ��ny�#�̙��f��)�9�$lg'$(�MC�,MǊN4Bzt������;}��k�u��1�n�~ڮ��eވW<P��}��WD�a��M��{ƴ�(�'R��ʲ��1O�i�Jh��L�G�Lm�-	���6@d�#�p*ư8�9r$����%ooo�K7��-=ou�h��!�4Q)-�1Z�52Ep���e�nT
C��V��$��%�;U/�p��7ބ���uBs%o�bC�-�%��꤭'��V��14�qӲ�Pu%��k�N��8]3��Y1�XZ{��$&Y_�=S-&���iD�Wj��zQ���@���_�В� @fH-�]A݋�2��%��ڗLǌr��PAkJA�����,���M�h����#N� Q*9ҚWvX�-��`��=4p�T����	�3�鏳a��-��j���w�D}Q���S�h�����d0Z�?E`�R�o�R��>�2m��:͸�6��Jh�f��e+,�+�ĚHR�*/hTf{AM[��C��c��!�A��D���$����ι����s:�Ս��%�Ky�oZ�5�Ϋh}��}��&���ű  !��
f����ޛO7Q�ر������ Y!�}V�ڿ�qS'O������R��WvR�%��T����h% qHڍo�/$�N��@�5���+2�W���L��ﬢ���m���u3y�_� {=��R���Q���~��ct���犰�fQ�0Y�O�)F�^T�7#$:�'W7�x>��2��g�Ym���x5��!Z٣����K���T��և�0�z)�ZRRU	�p�Ԃ"6�z�>.47�����>{��{U�Y��8�{0d�OC���f�of�Q�;,��F$r3��r��O�JvˬpB�[�o�k�?U8�`�գq x9��<���?+��_!�P�����Hs?<��w�<�t��O�+H�Ұ�ˊ$��1G>�i�~й 2�ѡ���بWc#s=1��<Zp�t���B�ZH��6U��yY�������,��§nB鉗rV=�J7��6�e��yTM��/��~��u���<ic���O3l"S�\��xZ8V������KxP�x�,��kP@~������E�3�_�d{ו}n��C���V��h<a���ۃ��U#��ю��J���S�;O��D�Œv�Ϝ
�w�z��S��[� �?Z�����rN?D����w]�GWVYD=���3�ե�A�h�;�I*�,#��fvz!�R�^���UG�6��>Tc�.A>x2p���+v��ƪn.$�aԇ�E�͋7n[h�wt4]���	w�υ�u���:8���ͨ�O&�j&��+E��?w���v���f���k�n�r���I�É�\ؐx*3�3�3��щ5�\��筠������5;��޴�uW������d�����҂I��ZpQ$����3S���Ek�1��8$@�!����>�;��L$0�q�Zu#��N���@�n'뀗>h�L�l�H�BR���C샖���"��;~Y邕���7Y�C��-�?�v�����U�_'Ae���Th�cKA���L��w�)��(�#���J���Ev���mk�;�/*1'N�������uEO��C���N�}��ޅ��Xg�IV��,���\ �q"�� �|a\K�~���bp�	�+�DyL�mv
eeژ���!&6ε��q�B�I�W��L�p�܆t'ۭ�?�EQw���҃`]��9\|Y��;=�(���Ow9�b��)���G��y��+�a]�g��V�Vo�}t�n���	�����B��,�4�41߮�a��ح:���;�x��'�6B\1�L��|
J�Q��N�;:���;*@���E��3p���$:Pv��� L�V*y�˩!�c��`�MAM�M���9z{���+aQ��_��\�$�}b@��t8h>p4�	�L\�@�Љ��&�v���g��ZH����L�T� FvM�!; Ƀqѵ7�����.�P����
#�3�����Gd�w�>��� l�Y�_U)�M�N� ���O ��aX*h2T�����8[���3%�&�Q�L�%�6���l~����s杚���ĵ�1��b�m����Χ2+�����;���C羸�M�Ķ��ךj�K�O�X�Q��ɞ�9+�_�B�6��3c� }�� w1c�@�ȗ��VK����֟���Bʂd�w��û�o|�'yL�`��$~���T9Y� a�3�1c9�XMQ��y��Ί*�b5�sgR7P��Q�cV�Zva
�*���T3�m��Ĉ��&$��q3���m5���Y���*SƑ|�s�^���p��x�:�e?�0cl��Y��R'b����0�s�rDT)���C�|:!�A��׽	�0���g��
!�ˮ�w�f�~օɫb�����ٕ��H���I�j+���~�B ]�71A
ޥi��	�?D�%{�a���	��h/o�\5Y�V�Y���-�3n6��%,*~�2H҂�?�
o�g�6+�_���>���Xr5���\���E����؊pX<F�]�K���^OI{G0];�����t/����cr\�����.���di�;��C'�rlj���'�LΖB�Vވ`#QYA���๜UpD
�������wA���8�%:݈���/�j?Ź�*��]��#��A#tu��%��a��+QJ�юt���	HU�4	/G n������;��$�Z�pkL?��b_p`%i�?�ަ���9,�G&���U����d�?���{-�5���SB$dWcx6���Ƕ�0O$���A������eF.�h牰XP��C�|�z��	W�����2o���?{���0*�������l!j"mn#q^\�ح��:�I=�� ح�Na��g>�Pw+����uqZؤ]=i,�b�m��n��_��.�o/c�r��d(n�_=���&PSk�Y��Y��b�<Oj;�'6�ِ�~f����[?�Z�>�� FA��tC9��6��.po����w���)�Rͯ�_7=���v�׶�9��,� 5�R|3�&���C�]pI�R:�90X�fs�2B��a�or���˔��QԌ�E��ۦƖBl9�:A��\���p��w(��T:M�(�g���	�~bh�	�.�*R�Q+�Բ�i=�0���v{=�)�4Y���1m��{ܢ���j/t����Y�k
��]�-B���5M.ȩh!K�{2�(R$TĹ�pJ񤡪۹�F��{�������["zS8���\���Jj%2m��p���o�^E�|Іm?N/�-�!��'� ��w,�r fC�����o�?�y|�Ť�2�#U��]���H�j1^&�6N��+d�
�d
�_ćNh�\!-wL����n�����?���:���JP��1�a��BUl�̻����6
S��ѧ�l��U�`�-% �����n�*�^^�g�|���@��B� q�~�DgA�A�J�bɬ��ֲT����y"#^�(.9"-�C�Pxy?���m�t\�P��]��o��79�9�B�1-�� �1Эy�&Wʙ���M�6�D�7h~�x)wv�G�G�o)R�-lb��A�hYI����$]�/}Y�0H���hT�nAAU:�����1@	@��Ӣ��K�Z��kt��=u�]�凲;�>}�9��x�LH��W5�y���@�1kw���A6V�/�!�\���~��<ޱ�ZX�%�7�e�ӽ�������H�Å��� ��n�ͭd}�~�^i=��TT��'^G#�C�Es�ܥ�(����R�J�y��a_8���]b�(�_YT8�m��j�Z��1"�gt�Jd^¶%,x�	K����*��1���j���,��M�
���&���i�O�m�GCP)&ĉ�5��-LN����Np�I^R���d�ʦ��p�@�Ҫ�	�H �(B��;R�d�G������p��g�{F�}�bż��
�1����mӳ����x��Z�r���eC #��K��)%�Y0%W�>dm����0gޘZ|��.l���g��>*�8�øƽ���+�Ƿ)�H�U�o-���i��=�cY&�t�@f&��P7�Zr��a��P�m�~�	�}����ԙ��{7Z��2��n�D���0��Wۍ����J<"Y.���D�J�U1�JT ��@��]C��v.A��K˶�����wlx��^�L~F(��U�I���ӛ!�\�T��yq��l?�&�x��7��
��-/' ω�3AHd�%�/0�$��3���3n�ܶYL0^L(V��['���"w����55���D�U}���Ł3WO������ƅɧ��8{��$��g}�ki���0:�X:�����¸�!��h^N���t��l�3'�ў9!�CK =�у$���U�t��z�f�q��-�����m�4���.k��2;b�� �j{�������(�Q9qm�L��O
�s���Y����<i����q���P����0#��a�p���P��D��MJ�G�A?�N�L���E��v��P�bu��q�#��^�jL>ьLP���C\k�I�������~~A��GC��}҈I֊�S����N^9�J"��G��|aC�2�s������U��ȜJ@��a���n�،�B�<0�	۱=K�c��|���(�F�k�ZK�^|
^q�@'EM��L;����ce缮��^J�
u�m�����U����K�b����<ũ��J��I��x���$H�_�н�?_)��c�F��?#,�k�f�Z���GaB�a�n����C߿~�'�Fz������عv�
`��	o��[m�e3���\�3O�/��ϻ���!x��V��)҇��� H:�a���N�th��i��-�#���W�9�~�D칃�C� �#J|L��A���3
l����V��r�Q͜�hn$�y���ȓ��A����K;��u�m"/Z:)���-��MJ���3��~�����otu��}�s�r�d�N#�K�y0���7�]�,:a���X�sn)YS�[�]�jl�W��=,�����qЮ���ߟ����V�o�W�OEN�&�*xS1]^����0/�?���ϒ���>����7��SA�|a�k�`�.��5À��*զ��/ʮ8=H��l�w�Hs�FI�Q=J�N�t�Q�LI߈����of��V#�
�%�Z��#��(�� �qs�`��}��v�
)Ly+��!����#vSq��v��"�m2H�]��?�r�js��l4��h�֕$��M��BD-]�?�8f����s���� ��/��Ü��	P�w<|8�W��XC���������=68�4�@������5O�w[��a�9�������pA��9(m��������ڎ��h��?�G��j�6�6�0��C�h��yoD�ܹ6ѻ���f<@��5���@z�fB_�ҥ ��+~��8E�R�|7.�s��Pի	VWr�f�B
L���&��C(��0�^�R���D�{�{���O�­��-cp�U8P��U�{���B��/]�w�m��X.�7�ߵ��E�W��!�*�՘�Eopf~�E��|`1�"��+Y��<�6s��/���@Ԥ�T�ȧ�MWmF�йϔ�i޷��g�s$�[�/
�M�`y�3���V�
�7*�l�u��h�`��&�$��
M����0aR7���rd�ʭ[��%d^(�;�k�`d>����B�n�M3��Z~��Y���tm������b�YoC�����x���;?��_m��j�M���6>f����p��b�0�-Z?�>�~&��^_��3&��{FJG����9��v���B�^�[s�=���&"~ƴ�^ pA��@9ޕٍs!�?�����Q�nmjsDp���E��J�F;K��a;!�r����d[�_n�;�Ѣ�j��݇ǑԜ���Dw�y\B�y
�ۃ�*��fA#mԢ�&]�Y3C��}n���s��e��7���f/t���MFQq��K-��
Uu9���D�G��P�V�]��x��(��'�D)�&�#��m�� A�y��pcG��<զ�,�&�������	fՖzz�>�g}��=�HSI����nb��6��օ�%G���T
��>{`���yVb&�a�J�勾��yNS��X/H�އ�.�o�S�ϭ�����(g�Yd�[�.�h�@��%��̯�q��~�P@�;]6R;0�����8��������co�+�U��E����}�9R�R��I����&��h���Y9�V�E�f|8��"��"3ʘ>�/���Qo9�jxn�ǼD���%@�g�g�Q�f}�hdC�1DC�bM�j~k�L�Q�S�4��MS��b���	�'9g��~ʨ�Ԟ�N�(��ui�#e��P'i,��+*�����\&FxI� b�2«R�뱭�@���ٕx��������$��"��S$hލoȑgxݎR���s�E�#��)9�I�v�^ܫ48��kW�o�� �[~S�yK�R�$e�.+���H��[���JL�z]�vl;���=��TSM
�����OG�o����2M���0��o�U7����t��B��(8eƋl��i~=�s祄����\��̢�{�$��&�DnH����\��A�z&ט;���c�48~�t��欘�q��^k���(��+;@���r�,�!S���٧��"ہ�P�,!��Z�ҏw���|�+����@�\v4��[�~&�Faſp��z������#!,�Dd$t�8wf:�zQ!^���V�V)�@���4ϐE�M� <y�l��Es��hS)�p�������cj�fӘ^�'�����b$smOU
����ѩ��JC����G��(�_���L�H�;"b�d�y�[Nb��V~�4�,��[���_W�|S� ����R�2��?m��>��5jgo�2���I*?��o�������L��ٜ�F�o[�R2�Unl�a��8��H�����d�}!��s��ޑ���vhQ#g�Ujeay�R����t���!'Lg��8�%��?-����aP��8��6��Op��#��QU�!�I΂�j�z��,�c�4\lٙ�
$Y���g�-)ݸ9�ۅ\����q8ٖk;z�b��h��K��.q-	�a�I��mB�f�(f������h�:���D�$"��!���X�F����׳$�iQ־;��ٴwl*5�+wd�i�C4�W�]�ލ�|��guR�<z���D���H:��I���]��e�%��y�\���J/�����"�Vy��U��|��̔���6Ý �Df�a".pj����uƧ�� ���Ϯ����n��M��8�/�"-�`v%F�ZƄ׊1��"�뫈:y�>�'�u��5/�x�Rm�qɇr����FV��d��z߽���I����2"��7spa�lw����,�`+P�.u�a)��� ��fU:�o�Ql���R�	�~-�3�|�"Z����</w ��'��M�.�>���੦5�����Ǆ�����F�Y���K�I�U� ��d���t��â�y�V��('�e; ��ƢU'u�S��	�"5�~$��S���tW�K�[�FT��OzC���k�ՈÏ|{�ǔ�:�B@K�o9��1kc.�"Q�d�=ܺ���f�%40��A��m�
�p�&�U��O���4��/*ƍS�����#M��rFR��Q�J~1�qm�|�{E���4�/���ߦ�4�����[��#�ӣi)c5΋�����ǩ�1�)ǠGB���ꨭ�
���7j ��eD�e�6�����m�j��o�|p���4�� ���}qѺ0�z�9Q\�q���)�d*;�I�����2�P�qh�E�j��ךj�e�ρP�����T���犵,��e<Q��W��b����
&� �E�.���8���}-F�2�Aj��w�L�x����D��$T���J�x�A$�&R��\8`�9]��i�0)6p���M?CO����\ՕR�E!f/L�����[Iڄn�9����q�@�,�����6� �Q�N�p9�J�|X)�fZ;=����(��v���X�����D����#���|7�ف�`",/'�����I�6�x��������j#g �@�� ]���e�����w��o��1��6��)r�rzBdA_K�;���~X���EJe���,�y���q>Ԅ�ӥk�z��i�5��:r �f�?�T
Ю�~�[�X�C��Y���煣�ܭ��qV�W��3�؜K�AԳ?<�́���ʩg��V_�$��_>vf�*�O(AC/�щ)(������N<����F��;6d3����<hr)̀ro�,��!�R҇:M�5�q-�I�(����n�����Q9}#A�dL �ۈ���$�a��SVr���!c&���"7���͇y�2�\��e�N�N�`�K��
�:�؆I� <q�@W�9��:>	���ӿr �`���c{v�J�7��uoy��/��,uES�:G��1��k1xC�<0��}W���Л���'jڱ������-�����Q�_����DP6%$��n��75���9C
Z���̷�~u�y�/	��ٽ�w�ˎ�#�a!���N�qS�+y�q�p�u8/�K�y��}U��S�ʱ�f�h�远�>[������h^��������n�A�O��0���1X�^+��4��X��EН]��~�	c��+`A$��;���l��F�!��O���
�����x���ѕϥzs�5�͋�D��O(��bT�^f����iv���R� �M�ة~[�I��P^{�P�T#�ۨ�R��ذ)�E�q�2/ő/ژ�#K��*��)4��\�A��8�kЦ����J�Y�0��]��x�s��?Źs��L;��R+�$7��$��]�MLfg*�d�����p������Pk�C�G��+YG�ӄi�ŋ\��������O��^\#����]WD��C� nY�sGnP�?U$=J�l�B�dw�lXZ_&�ؐ��K�Af�9Y����,��<\,�ߍA�$�x�H2��w[E��Х���ADn`�z��`��d���2R��AFJ/$�I�l��c�m���d�Pu�Y(�>��O��=����� ���&w�=�( X��&�a8�F�X��x�'-���J�G�ME�LM��#s�𵾴�5(�{Q|��ݮ��z��w&�X�;.P�r�t0w�[�[{@����R�l��{=#d�}O1�e$�.��N�ͯ�|? o�����htӭ��|;�1�|�.���*p��^�r��&=!p�S�?6F�f[I:�;�	@WFq�k�AW�,x�A��F������d��\H�8��2�r ��m�C�q[��{�hp��7z���%��U����#.-)�q�Is������R]I&ʙ�wS�"G|z��HSi�[!����A��3��r�N��R[�k� �[�������<S1�-k SKv'A�Q�Ə�Y2��0��w6����>�k8���Y�81_֫h�R���Fq����$�>˗1 �pz�`TaE�����i��l�D�Ȫ��O.9���*�x6g�{����}~���.�����b=�z7��Y�p oz���S��d�Qk@��n괡�{p�!7C���'�6��;�o�^����F�X�dK`�F��[a�H �:���-�j:,m��l�yzI��w��4��j�WuaI�������`�ؐ?��iF�q
�	Uʣ_T�$x<�纽��6�X�����q���Ɖ���{�	�������1�|d�lp+���#��CLj�X����#Ι�k�f[�k��d�gr|��W�t��0����pi�����w�v��q?���hU^
2C"���a|4%���zV�kY�pp{�W��_�b)��F$� ��˃�i��� ��j��ZP��v$穡�+P��0�5a_��
�pd��;��)78U�����F
M+�ٱ�ؾk^�Ϗ��RvQ<e���C���s|zƒ0dDI}O9�0�<C�aZ�=�S�4�HK;%0�_��ben[1��+�o�hC��1�������|�Q�+@����.�Q�I��ipLF����X%g���U�>��q�.��)�O�l���jD�@�P�g��7�/�y���6��9���5d�m���*Z������|�	�����<���q�C{k<T���fw���Fr|�G��.�H���Y�z���0?��~�i���iBҬ��6 ��bȎ�����S�D
ʼ��=�H�`:q�"u_Ф��BMJ��L6Lq��8YĞ��KZ߄-�$���X�O�W�8�MK�&_��r�le�h��VL���d�����ӟi�Ǧ>�D���H�|��~B��vQ`�t��_���u
�^��g��<2�	�±$��H����Y޽�h(H��X�Hg6�XC��v��[:�.��5'��i�#�_=�-��9n�P=(f��5�	]� c���vk&���/��;�J�>�ޔ�����~�^:���Ј��	��9d6��!���5���r�vk�d��+.�c-@ĉ��)ʰ�j����/ܝ�{��hгF����S��&HE� Y�S�8�<n�r��ˌw��3�|�a\�~�?t�w���3��"W\�%���qHB4�?O�U�2p�t���F�xgڥ�� �m7D$���ЪX���٤��-�ȸ`*���r�9-����^i0E�\mp>��j����^A���oB�)j�=�I�?~i�Z6؟�����vLuၸ�#��DQ���ܱ�R)���,��A&�,�8�FGmܴ١� ���=W�m��t��D	�g��Ul�<&FtAA�Mv7�S=�t�����caf�Qpk���-Pd�*:#�ǹD_U����[NHKn%�n	�w����Q_�\!��-�"Y�^���#�s2ݿ��$h٨]�[���">��dG����)U�� ��Ұ^��j��*A�O@W@���? '�k�]T�t�,3*�M�\?
b�k�(8����ֵl��9i��Q���&�f�K��b����+��j�%�s�8qto�������d�#�+`̭�'H�H�k_��dv� Gk��vJ������u;��U�/�o,�O�C
 �TT)�v�B�HwI��@40��P�c&�>����r� ~f��̙��ಽ��B�����p�!(�^��3p�"����.��X�tA�fT2�G�<���R���������� fn�5Qڮ��3L�4?P�u�r>�p��D[�0 ��o�"����>u���g����k�3|9!����1SxU��:��a�,/+�0"]��}�j�G���wv�ן0�V��Ylf�"!�݃?�G��d��������2v�6��j��H~ʚ���($�'*g������*�P�	�A�3��ǛyW����Q�S���e�@a��RW$��Yz�H#����^����kN��b5DK�38+��RZ+��6��ۯ�Ry�b��Ӱ�����GE�L�4{����ᙙ=p�X=\+��%�=3^���%d'�G��̄��*��=�J����>�WwV\�̿���A!Ъ)���)��2��Yѯ���;� ��
<�_s�	�쏻h^+����zs��Վ��} Ìi�������t�1eV��A���ՊE��m��L�~��F�h}X���ʃ4Q�@�S�@��л5��l�<uB�IhM�)i�?9�q���X�k�7�Ho>�K:gEq�c�\&�Ȥz�f�Xf��,.6�B�&gW�*v�-*����H��_q_�o{�V;g��ΗPTBۏ�U���8���5������W2Ř����ŵ*�2[���k�_�@�+��=���[�������BT�O]����� $o�o	,dϞO:q^_z�@��<���`�] eP~��O��62	�5N�:#��0��p	��F���(J����--[4=$]X��N�<�!u�T�T"�A�@�H�Hi���q0l2���
�p;�QR:]oi,�:�}�,,5�(�f�I�)F����/��+W(�훤Щ+�GKB�1�J��͍�lC��x����6S�}��k��@��/Q6��OPL���V���T�5)�l�7߭j*�!�mM����Lj���iǌ�z����.�7y�򉛎��+�Q��������l4MѨJ��%�w�W��
�ْQ؞Bӟ���* h+.g�ׇ�z�>|&z�S����,{d�p�K����zg�|Z�'V�n/;IVpRJx�QLV��K���&�q���:2	�3W����ky�sJy�U�	!�(�������?VФ�I(�ٛ�B:��}u]^<GOa����\�8x:�*0,��b�����v�)�����lH��D���r$�����Gl�
-t��j�Ű��v���*e:�q���Q�W�7T�g����f����u�Z,�H0�I���j )G�R�O��6$���"�9�:Z�/ܖ�'Sk���yV��Rĝ@��[�5���.QcE��N�wM�9�Z*�~���uzj�yK��潤�}W(O����������e�#5�2%X��x>�Y���&(䘵W9!��;�ty�5SSö`~�ǆ&:��I�l{8�ȼ\�.8Tm#>Ԏ�c�][aW8���=Y1t���U�!z�%=&�uI�~��.�L�!vg��������ծ���團����9=*���w+N���N�Q�M�rq��S���I򣆴�V'���@��U��w���][xH��v��njF�k/��/u��ĸ�<dŇb�K�%s?Ht��X���������)��^�@�,~кqG��rF�?�C%<���(G2�@Ι9�|;���4������|4c�@懰��h /�3P�NnVQ`gY2Iu+�����4�-�!�[�$�嬊������n�]	�ݑ��@�;���~O�~\��x&/*�����Lf��xA�+=�����r�:d'��x㴔����fꞍϵ�n_�̫�0�i4�=`�0�'��;�\|����^�-������h̕���������t�Џqh�m�'B��1���I��*s����f0ʒOcE��W)%A��R��|1���GN���� �z�� �۫�w��-(G��F,[��>J���nS^�����)
�^v��+q���x����H�+lտ�/��z.����t3�3y-#����?W���p�U��ߔ�� =7�n���:��3�P�#���Q|_�����Ԙ�&2���b���}ҸcucSȎ����8⊊��v�����`�@'���0[�Y����2X��k
��ba+����h*c�ʚ@NG�7�gZP�Ӡ�3���d�#�� �w,�I�zO����½ϔ��h"^gZ�f�.��SU�9P&Z	rDѐ�Bu��۔0���MeҋC~�"z�K�q� �@�zcθ�d�����j�8�N�0A�㫵��IT44��$9�q���b��U�x7��94P7� ��@TE	�����t�����K�;\b���,�03��i �a�9��~+�>XU�����մ��[�n3����}\`�����q5"�FP=26g����;�|�/29o$5lqI��{��q�m��މ�P"b��L�>�;�K�n� x�e��� ��l��\�&��E(R<���)
��)��]�f��-����X�^���|8!�N�м��G\(��hZ���*�����zl�wfT�D$T;*=Y��ĴW��؏3��*�f5�L�����@�D��(	�^���Uy]��z
+.�qn���[TQ�L��'a�ot�t�nb� ~�?�.v�g��r۳f0R>��\��$�=���n`I~ڬ��Wj����CtT�KDz�L/��#,裠���Ш�0��jE�=tes�?*\KT����n�-e�#D�����B��� ?����b\h��*Q��E�/"�wsCM	i��cXecQ�@z6�[�}G O�t9�`�&��l�����w?�n��Y����K���kJ�i��Lc{��+�t�Kt�H�p��e�b�!wS$��{�8��c�mw��J�T�}KA��"�&���PqωJ_R�6����\���p�dfU� C�//H�ᾺϽ�����X��I�bbJG��$�uur{��+�Yc�Wdf���[�RuUQC�N��Z���v*x����?i�E��z��뗢Xv��k�/�6��7X�O�I�����D6����������6�ݩ��
*����Vz��)w���-�0�>���6Tv���xlC�N��nf���S�ҥb��3%^�S/��;���T��R!Zvۓ�����&�{��F"�Uu��2څ4�+��g���D�,�'��aQ�q��1�"�I45�����H��Yo�Ϭ��"�f�@�?f{0dcmo=�h�������WE6��L���y§K�0~4���o�^����)���N�\��RjU�YI���<16�Ml��
��tHQ����l\��A�Է3(`��
TZ���:�5�[��u�L�<7��UhYO�kBem%� ���	n�"1�!�G
x��)������@��i�����-ӷ`Ψ�}������#��n���b�'C(��$��OoҭKa��R��5�,�(�u�����c���}���{D6���cU��V
�5��E���B�\��_VM�<��nP;�2�ҬWR�ދ��+�&�ٝ@�q�N�,EJ$�9��c��P�GJ��D��c���E�(<ZKNRmԑqs�j��a����q�@��u/~�T:2q�W�]?�&��m��_]B����5�^��ƀ쟞r���`�3�6�S��և��{�<4�F�|�Cb2Dc�a�8��{#�5��m�� �0�i�)�O}��h���Ie�h��s��y���uoH_����2��:Um��)o�ʀ���æ	ho�+7���n~Q� <M(hد�_1�GZ��)H��f�"`����@�Z�*�8��������鶮�(���,�;=%If�T�������XQ�Ε�U���VkU���Y�̰�hR9Z�<ؿ�q��^&͈��
�cO_H@�'8�!T�J�jUS��D7�.c��A3�2�/W�(|ke�O�ăxqp�n��'� 9�.�'�O���W���4t�����u��[%����M�@E����Q 	;+��vj(Fzi��(�\��]�.Rz�2�e�8��l�B,`�TgРK�R��"Kp�73��� �&M�>�椘�5��&�!u�[o����ǧ���XSe�sn+�Gm�@���7�.�-�[���F�:�k�U'>���8��U�t��7�M	�B�5,S�y�8O��!h1�e�f��̳=T��CD`�'�.�\ߠѣu��v�	�cm�p-vD��[�!0?�i�����90M���*@@����6��W̯�)2w�b���I���I#\�ʧ7w�˵k7KUo�t�qT��L�7&�Uǚ�'	�@]�՗������1�J��i�a�5�t��^)�Qb��Bc�˶u,i�s���o,2�[�ua�I����M������l�v�P�
~!���نB����R#�G:8�[Z�٦Ub�(��d��-�/ύ�_��~�R$�,K��e,N��*"ϲ��	6����������{L��{�Nn~�ui���K]&^0�3fI�qeQ������c/�]���C{��M)�Qǒ��U��/^ǚ���Bg��ߐ��q�D��w{w���ch��	���w��כՔQoH̳Fc��LB\(^(��{�����?�x|�� �!(������,���PH���-$U$ꧺ��Ϊ��z�g�`F�L.x���;�fi�?�
���
.}R��g��.J���kvڿV����&��?�RD��~�!3�g�#���Q/��n�t,$��6҇d��Z� �.�<hH���+P.�*�H	�ZPJ���:4S��S�Y����6=�ZG��B7lOK���2���`8q���k�p�@�&��F����1��+_{@��n�ϘC�͙�oHu�wz���׭�=?�U�=(bFs[�y*��V�E� G����`�o�b����,���sh��(/�4��*%�����[�0+dʜ�P,T��hA���Z$�]�#��eM��>/Ȋm�qܢq�sb��nATq�(R+(A��D.��:t]�Y�o7��W��G1,���|� :��3����ܙ��>3�w�Y��̑��,��D�Fl�6([�� 2�e��L!�4����0~��!�s(�j������N�:~wd���	H�Ƀ�٠�~�|о��ɞ�t(��[�@0F��t�#�./'BX5	y��QD�K)�V�N'HzR1=�:᝼����қO�`*N�\��.��%h�8�W��O�0�x1��*�?�&�1M��*rr�ž]��K�:���R@��l���s1��7s���MI��͖���j#���v[�I��k�J�|l�]��_m�"�G��A�A#��~��e�Vp��n�����r��ʷ��?�ډT���>��3�/C�z���7����}1#Q���׵AO`��dk�	R��S�����P��#5�}��+����������l���cG󓢉ּ'��Q@JM�孶^�:=�Ĵ���Q�jtщR}�{��|����#+=�.��2��k�\
��	+��u�Uj����ܒ�;�*v@���z���M����
���s� 跴%r�<��Eh���ܷ�xJ_tBJ�תz�F�LX�(����rY��0�٤�2�/:_��.���ɢr�fq
G�;|-P4�% �!�{�O�KQf�"�dژ�z��og *�	���$Ξ���g�y�)�/��7�R4+23�S,�,��l�y�D^�����Y�ʨ�="%�������UԚiZ�Y(�8ے�5M��ۃ&=_�֦�o����*�Y��-����۱W��-x�4�;���KB�'�K�1Q4ʺ�e�b��TFeGz�k�K��2�RCy�BJ*Щ��a��S���o|Ő������e�į��8H�P�Lz�19{�]�m P`컣�e�"�p֊��ji%UD.�����
q^�VUɜ����-hӾ��Gl,`FW�^�u�9��k�/(���LJ�sm mA7�?nуN˚�F#��p��$n7� Iw�(�d�'�M�����9��+	�?:c;pP�B'ŝs��KC��kv�������j���y����m���ܳ���f�O�"ԐʽSr�v�!i�)eCHx©w�`��3�����@��n+낮�:+����Y@���`є�>�:��Ne��o�ez��v�0/0�ur�
v��"�Q+��R2KV�O��Xթp<��^	f�Y�cBX����I�G2�VSò�[��Ls*X�C�͠�E1e|�J!o|�2�
A��Gr()?|�t�̀1M�mD[(	g����vy���E
�[��ͱ�r�/�{��6↑A/~���� ��xYi�y��[v�]��,ȇ��7����l 7W�Z��Vji�B�S��61���/�4��^�/�ڋ�K+�j��#m�&�B���䎿G��h��pY�7鲫x�>2©r�t\��>�s�n��g�0��������!Aё��L���ܱߥJwR���7����(#'ȅ���ԢO'u��d˔�èL��?�s�x���%�?S	��v�B{9�7wi7�1:vd����͒5�wU���8��C�
)�����.Vu� ��9���&�^o3���=��26��1[��gw[�v5�9�� ���Ɂ@@��~�_�l�ޜ`�$�1�a/Ы|���cD�q��J�גk����p�K�Ӫ���Z�=����8��V{ga>� ȋ8Ӵ��g̍� �ヲm�J�(I��ۄ��kO���²�sU��tp;��9��M��UGvk�xsz��K���N�����:E���X�a��E'�[e,F�U��_
��d3Q�>���PI�	!>bd얅N�S~��k�Ye�-���ɱo��q�P�'����F�#Pq����j�ů���<E�u2u�}�g{�3��zy&���{�^��-�ץ/��l!��*�֢�k�w�L5aqO)րa�UtٙJ��%0�5��~-�A�0�6����q#�YR�x�EL6���ݮ|.V߭�^ ���A�d-�\�Ϙ����wU�J/��k/���a�EJ:�'2J^/�ܔ�b����ϸ�R�`EE7n��`���0�J� v.b��S8C�vN���L����z	�٩�{�����(��Q��{��;!X۶��A�0�4$��B^0���-�i�j�F�O�,��8Z��ً3�O8��y�f�77H�Q����C:�$�,��˨4;V5r��.%o\-�v]B��P�޷��WA~��q�t������o:_H&����D:��X�My����F�$����|L+��.!�a,>�|���������A��K\u'٧.v긐�8!����n����`�T���{>�oL{C��޾���O����j?��-2�hÉK>�=G�%��R'C]qƧW��N9�3���w��t��(�[��� ���=aa�+5괒�I_q�7k�JT���T�+�=^���N��v�j���2�|ׅ3٣L^�j�ͨLW|)H+&�/��U�-�ԧ2�yXU��J��;�?᭻���F
i)|������/	X�h"Z4^~�d��x�zgIxcu���c�"�d�ފ�ߛI����;Օ�������TՓa�q�M�ʒ�n� ,f���H�Ů��J^1_Y��M��a�@z�/)1_�������,��%0.�w%���Ze:&�
��
2�%1��V��g+]��.N-z�7�77���ĆO^"�ߺ��,pX ^����ps�x��]ْ<?��re���\�L !|^��R�ǹ���7t��/����"��Sm4Y����"=PzNj�
�:��3p��LŠ�i��<Cb��P�>oގ�޽�c�<�e?g��>��&���fw���^$�8�P�:*n1�#a5�Y+�фg)+q�r�����0�����,\ �a9�#49�|�ا�`�Ηd�p��.��z��ދq��z���K^e��g�~̐�c�����k�f8�>~e��R[V���Bd���+�}zty��S�@�G��~�:C��{�kAm��Do�N�hm�m��daC��=A��� �O
����+�R���c��XE���ʞO�Y�Lb��k���L� 'e�����^�>D&n09�Tz�o���|���v��]�q�{
��8ۂ.0��tMj5j��x�i۴�0Z�W�_NC�R�S��"�~:�N�=�eV���U{��r@U�P���� S��Ir{Dr}�	�S��n�v��ݐ��������|^q��ಥ��|O�����D/�n���B�=�[�o��? ,��n��H��'r9V�cD�I1༩����i�H``�	�t��b�]���*���"��R�m �\��􅽨�P��6Fl�"�M0���__����Azlf/{5�^�3�����,�'�%���Y@r�D�1"u�RLs"M��{���**�FX@��a�����J�Ӓ�T�J#����&V�I�&�}�������l?H�#���l]+���pH�h��u�^�����ۯk����A�8lu����o�q�L�Tq\tX?x���� T�TZ�@J�xb i�^
���=�9c����J:JC�W��Df��gf�í���a[��_� ۸�Ǚ����L�]�;�W�BqS�k��S�~.�>r�Y�0e��� �=ܷ-;iv��p�j�+�2+t�K!3,"�AS/�9[-i�0ן�ǻ����&�)q�U"Ac�U"� ,2̾ۮ�x1�"����X�b��(,��AN�o��]�[�@��DG�I�FB"�>x�[�_���F���ϑ��R��TQi�i��	��'��i�`,���}
�ĸ�)@+E���������c֭�:�ј3 Bj���<d��\��^��)��M���M�"�0���U�5C�E�]a�n�E:r�U��s�)���0]��!Np! �$u"Q�� d�"�2�O�R����^|��D�[w���ȓ���H�
��5���A�"~�����V��j�{>�e�����r��f�ЖRTp�(��?�KiWpd���)���S%��U�4�u�(�T��GL���M�����	��b�<tc����-�*��I|��H�WzF5&fa$`.�9xײD����6�g2M>N@c��tw�
Z]�A���
# �n�chՄկd�R1�crE���\cj��s�����*|ɓI��IG#��!l#�ZU�W;� ���5i�N�t��ߊDu�D�f'���T�:;���u����cs2`��*鶾�E�����gz���0����ruN�D��b�4�&Ε��](dA�g����[bvx0ɁA�A�th�%������uW�u���uQ��$�@��zlMN�9�ם<gD�̵73b��!oh��Z����ν���B�џΈۃ9���I�n���6RL�og��/t��z��{ao�?���P�w���_�4 O:q$꽹�:�ȖV�8)�({7��b��O�Dfw���y�T7�����K��ÔJ��I���W���ˬ̄̇"=��r06
x/\����nSú�M�
�N��yK����%�ETv���x�Nn5eo/[��u��uql���iTTG�z`�����R9I9G;"��x�z���ȂSנ̃v�!�OcΘ���ڡ��,�L�g��Ή�g�y�O\�Z	2��+�жB���F��7�O�$��*j�\׼��O�1֒��Ͱ�����*`��A='K;���t_~2��h���cbp��[$ 	�g�l6��1��j�Ь�s��]U��XE'��@�ԛ��T�&~%�z�+"�B�X��������ʊ`��s�T��MfO	o	��n;�7Z���*��q�����;�H�O�sx\��O9(��`��UR*�r*�7�Y0#���$�G���R�H*c���1��X�3�/�I�A�9���Qݕ�`Nwq�u��:���a�� r3Kj&Dε��qU��gɂ�c���yѽO�� �Yo�����~��[I�]����\ 6�U�R/��W�'�/��e��_�$,�'t3��X�eL�q��R��s��Z���0`��>��f�>l��V���Jd2.b��l(��&��e�`C�C�I1H�R/��k�+����6������P5�C�������W�Z�X�[tܕ���+)��0�au+݉�����e($6nm����ڜUL^�U<=l���p����� ����"�[Z��O�5E*LhY:�gò���Ҋ����}��k6���i��fa�ˬ��s::h7F��&�F�,�����t�I�m��GKm�o.w���0���^8��8S�����@�iIVH�bc�����k�pk`N7����l�;M����$y!�F� ��ob]*O?�Vg��N92y �:G�
E�0��r�IF���vT�^�_�xVk�