��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��,�y�}�ǰ�=4d�H���`I"��W�`r���T:tB�T4D�m�)�	1��I�t��
��8(�8t>s)ו�."[�漆���]�~�]��;�O(1#5�-� 偙O��QZ��~rL'�x[�i,mׇp���O�I43��4d�,�H�����SN��d���3���r��m���̨T�I;uj2Y� Er�*p�Q$Gm���p�V�`�2^���,hz�<p��l�Bxt�5��s��\yq���#�@W���f:m��T�	,*�񞭋����_��㧋l�	�\�:��uGd��PǷ��N�I��_����Tuv� ���us�(H�~�{2H�:Zor�Q	#%�3ˠ!��iS��95�,?�.���/�F�i{#���Tp5����Ҥ0{%���2vpn���X�����@l����3dc�ק�3	�Ed&3�ZN O���z��s�yxӡt��v*}ԫy nj#��lc��m戭k[��5)�A#�����8�!�]�Z�s�M���t��w�!��'ÒE�rv��Ϝ�c@<U��\tq+��&|�&X1)C�����r�A~��B�&�����s�:n{p��͠R�X⺂L^��R����c���f��J^?��ܣR�O 1�rV���:��T�4���AD����˩�F�w��)Dm�O�b,�a���1$��c��7t[i2>�ޔ0,S���󧇳Ϟ�ᒨ�-��}�!6��Jyv�醊�^_�(�H�(y^����o#����X��3-�k\8�M�T�"`R�DF6ȕ� �,5�;Ҭ C�k���1\������k�t־9�}���� ���QHF��"��t�9 ?��{E_�7��!����](�S��0�q��w�9��=�i]�1�GʦȪc�W�XC�|�$��}q�6����zf(����լml�dz������*�eLD�*�,�m�]ہ6����D�Gw� �g��' A��)�m���b��ӎ���o�6ūvO��=�W�������}��	����z
��z�&�P�K#�^Qץ�_������&�)�ٺ�u#uD�	' �/|�qf�M&P)�tL�x�?�u�����ҽ�����*c"q/�\��YDl2n֢�vtX��Q������ǰ�6K�gVL��ο��Q�������-�˚e��"gb�_� L01�D��ثU�8-��Nw�@�$[�>V,���6�����=����{>G6��v�����φ+Y��	�d�A��b<�)��Gp���k�(�vWu����!5�i�;�x�60V`	��r�&������#sy��F�$�('N�w����,��	�+�H�ڰ2�1FÍ�XI�F�w/��i�Tt8"52�� �	��������tU�����O���-knr��ˇ��@yP�Y�a��]��R��e�%� ��[,-��W����g�Ւc�祑/a��l�h[iHk�ǵ��=ڎe%<����E�j��������m�(;[]�����x*R�ˉ4W~�T��Ȉ8�B1�� ��#�Oc�/or�q���Ȱ�f�'�~��Q̐�;L@x�]qK0�{�ٿg�b��	j6�Pd\Ʒ�?�i;,B��,{�㬹�ލ�\�a8-X	��{aW��h:>k'c����m����i��0��yn,�m�3�	�����, Á�J�/d�u `��(h�O)M���m��W���pA굯[���q끽�/��E��4-������״2tç�8��g�u�b}D�o�Z����z:��Ф@����f,��U<�yt�Wp3��Q�-a����o��]�i��ˁq] ������-�����M�c��8�ύ?��0�ٌ�w*Y`�뫂�OU�0��8���M�=�Ҹ������aV�>����'2��L�՚� ���
�ޒ�K)	*�#`K���L8P&� ��������u&�}G[>:�K�\��gg05�abr)5ob	�nW�����\�:M�WT	p����%���c	��Dp�[���4@m�W����!�!F�&w=r�Cv|�b���Ux�]�q1c�����k�C�x��g^ж�k-���A���I+/�
i3�W��cN}���>+�q]�6 �N�Z����ꈻuTQU�j�=�
����ָ��p5&�xV	�|�1M��lx#	��;Y�o"���K�'~�@�L�_�^�8��<w�i�-�sDq.����A W���'���{����$��ڠD?FV�T'�p�Z۽=��r� �3�ۥT�N�:~����D�mcr>?����RQ�-����Hr�8�Yzq�,r���Z��Q�[�>�M'�w���0x) ��i�}��HN�ue�	b��F��5�
{�H��Ӱ ~v�ՈO^W)̞�/s��5kYh�"�YeV�_r�m�j���+�k	&��H��%6�(=	�����:��#�[��`�͐��ohW3c9	�~j�4����}R��˃�'2�>��Fl�f	���r�ޣ����KM����rAq:W	�(К�T����m�^�FG<w�*�����Z������Y7�f�����S��+Ƶ���pcB�6�ScD���0+�Ԕr牰Y���@���.��L(����\��d�Yp$z��0X.�}�3�>c:h�S�ؠ�:�+;d�*D�G'V�4��őm��\d'��vMS����
��P*GX��A�,?���;�I���T��鯎�t�/G��!�gA�����>�Tj�Yv%1���� ��>����!�S����j$s�������z�~aN�̨y��O7N�_9j����~;i����Z���-��v���c���x�T�iߑ����i㴗���ƛa
���1˼����� h5\}5^���@St]H�$��0��t��O�:��[)�m�V%�"���L��_���d-��l���.lϊ�����O\��W��-)M%mpU���<5����P&�	g�~���&tk�:f�����0��U�^�l�I7�3�������~\�{؏<6hS���u�lmr�/�C����@2� +v��/fV�ۺ�6V��?�X~�՞]T*����������h��n��e���XO�=��+�>�<U}$��\U|�ۀ7��ƒ�_Z۫Ĭ%���.�d���>�h`�����R�H��2�L:��������n.����!���Lp��3:�H�u��zFW �y����4��?��N�U�MTY��qo�bǎ��d����9�<�[%�W�M�\���F	�j$��E֒��.�_�������Q3䰁�	�D���:�
�k��u�Hr�+��s�ndS�⋢�2���?���2;<���X����K,lƁ����scltW��u���H�?��OtZ(x�v����`�ևVR(��Ã�^,.TlZ�W���G8zL�{�Ʒ�*���:7m�oUǻ�wZ��:�w��iY
nݹ=�v	�K�g�ا�ˈJ�O����jѠ�VЩǍ2�9«d�3}ܱ���.�ί����(�6�and����H�}Y���g���Au���1��Z>��~P��T9�AY*�SM�94��S�/$���;��2�J���5vs��Xd�v�n�ۥ�h%���kyՐ�Թ��?�zUu��';&�bڐk�Z[�-to$��-�v˺Ʋe�ڤd��%B�X���Y�nC�y���>er~zk87�z����{@�q�6�کՋ��4R���d����ړ��j�̵�1�P����:}�+X4R������ x��\����a#����
�)aMms�j[��˟�O/$4����8�x����T>xt���m�K�״���"��ww�A~���@|,����J����L�����Ƹ5z��;�>��e
}dSu'�����$�3zI� �g�M1�s8��~HV�_��b�j��{�J*��fVN�"�R�C&8AR�-;85���!��gC���|T����S�t�ڧ����߮��m"R��F��.��<��Hh�0h�z�CM����6���^J	�T�-j�3�P<2(�Q5"��
i�y@��W����X|�g��9^�)��=>
w�]a�Y�,��M����t�+3n?��! "Jp���[6):�-�%9���q�<��O� �T'3��xB�f��w~ީ'�k��q!��<G���:7��vU�L���S�'��Ͼ�t(�C��.L�Tְ)�0ǤES_%�l7�;��'�e2\97ȏ]��� �Z��S�^���A�E���A���c@����_�A�ڴO���]�Jq�n��-���)�u�|9�,{����7�euJT�~���6��4�9J`AnRzW�˚U�7�QN��g���WV�Vd˭벆MS�:C��Ь���Pgg��^>�n��������[��,��Q+%7��}/_��t"�{�x��ֵ���I�&�89��1����UK�E�'��G,c�A*6+����������<�Ed�l���Jh�>��fN�-z�:��l���4@Lֲy��7��}t�`�֨a3J�Y/��0�	��CJ�������i�vWƪ�[C����ܸ�o
�����Ujȇ��H2]�X�˰R�N�]��y��E���
=�vA �צ΃���7�%|� ����������Dxk���� 5�b��D�j0C
*>z��O}%ҹ_w�h�c��$�*�P+2�:�O,e��ɡ�S���7��m�1���G0zJ5'��Fv]���y����~Q��� m�,ј�!jw�=ٛ��fDٿH|��;���;$�1��$s�"�%{W��<�q���$I}Ň� ��q��_1�+�O��z�=Lkm�d��C\J���9!�:�\g�U2�>�	�Yxd��Z������q2���b�ǖ��_��R�0�!��Y"Fԉ��k�L�4�T�m8�9vx�3�
��ZG�T�[�{=��fb&�Q=?���G�n#ᛥ��j��4̜K)���������oJ�%m��)o�d2�m	��X�E��w�`y���H�gzGJ�u+�I�k8-�m|[�;v$v��N���~ ��W�Vt$<�uϻzqO���H�����L�F*>W���j3$e�\T1��RD�E�0�J�<�x�.b�2
D&;L"[�Viʟ���g�u��V��֌HՑ�N/�gK6��g����^pn��/^e�=���<�]ˉ]�R�y�Y �l��N�>F���v�����'�Wuzl��7G�/�5�`R��7B�~���6�:]s���L�R'�	5�h�/a��ZD(��\ع����<tMt&�+��e#��J8�"�/tP�5�!�]�����ցY�}�[ ������K��̀�Է�<��c��1�Ը䵉}��]MDˊ��"4
$��h����CU|u����rA� �_��M^9���k�z���9g ��9:	V��,V��e"�;O� E�j/eV�E����w���K�-�`d ��X���y���W,��p�g�»K2������!��-� �d�����p��F���&t�o��t�*�#�@���`KXK�TJ�kn�|���WDC��A|��#&G��5˂TEu4%�t�9��#�Uk����`L�i�<I�10��mKb�x3v���Q�\�QJ��G�@��T���2�Oi�)�ۂ&o��
d��<�y��̻��@Y��g��Y���½��Vbz������4<@�"�"���6[ɞ��tw��Z�N!C�isg(�����֙2��d7��[�Ò&���㐂+���"�f5{r�($����j�5^<س�������-1!ȰY�/��Zmmh�M�Xx���xo�E/�fӫ4,�"L�BG��"����ׂpØ�9���A�j!��M�JV`�ͣ�g�v�*ta�ʖUb�z9� ��lH�Npa�y*?� ��Y�p���#*�,^�B!@�M27{~��#�8eS .:�_�