��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��,�y�}�ǰ�=4d�H���`I"��W�`r���T:tB�T4D�m�)�	1��I�t��
��8(�8t>s)ו�."[�漆���]�~�]��;�O(1#5�-� 偙O��QZ��~rL'�x[�i,mׇp���O�I43��4d�,�H�����SN��d���3���r��m���̨T�I;uj2Y� Er�*p�Q$Gm���p�V�`�2^���,hz�<p��l�Bxt�5��s��\yq���#�@W���f:m��T�	,*�񞭋����_��㧋l�	�\�:��uGd��PǷ��N�I��_����Tuv� ���us�(H�~�{2H�:Zor�Q	#%�3ˠ!��iS��95�,?�.���/�F�i{#���Tp5����Ҥ0{%���2vpn���X�����@l����3dc�ק�3	�Ed&3�ZN O���z��s�yxӡt��v*}ԫy nj#��lc��m戭k[��5)�A#�����8�!�]�Z�s�M���t��w�!��'ÒE�rv��Ϝ�c@<U��\tq+��&|�&X1)C�����r�A~��B�&�����s�:n{p��͠R�X⺂L^��R����c���f��J^?��ܣR�O 1�rV���:��T�4���AD����˩�F�w��)Dm�O�b,�a���1$��c��7t[i2>�ޔ0,S���󧇳Ϟ�ᒨ�-��}�!6��Jyv�醊�^_�(�H�(y^����o#����X��3-�k\8�M�T�"`R�DF6ȕ� �,5�;Ҭ C�k���1\������k�t־9�}���� ���QHF��"��t�9 ?��{E_�7��!����](�S��0�q��w�9��=�i]�1�GʦȪc�W�XC�|�$��}q�6����zf(����լml�dz������*�eLD�*�,�m�]ہ6����D�Gw� �g��' A��)�m���b��ӎ���o�6ūvO��=�W�������}��	����z
��z�&�P�K#�^Qץ�_������&�)�ٺ�O�? ~��@`������M�����@��������$	�(��%���>�*������5�m@���E#_���k(I����2"�h���_�]SNv�@gԁ�5�%�����O�1`?@�v]?�z�%��8�;�e���o���(d���0{�t2��ϙ�!Nl!߹�oU��/�0�c"Ӄ��_{z�}�9^&� u�]1w��砥�E�H"�F�}�8�`�%w��Zy��5	'���.n!�4@���1�ԤXy�rF��}	#��U�nz��Ź����$w�+��.O�UL%�Ж�kVEW�q,����%�M���2������4�9Y��WlYA�*O��ުF�A���J'��޵�{ց:C��\��<?h�^ �J�:��7:��e�.9b";)Il�o=�j�*��+��Ч���$�q���{M�^�u[e;wd/\��z���z���N�"VAw��f��D!�b�0\J� �_c�(�Qi
;�=�����;7a�a��a�	�ρz��4ˌK$`l�'{O�Ao�cV�Je�q'�4^�4���ߥ9E7Ly�$�M�ro�j��b����Y`h$+���u�j7�]���(�'�J+r�־pvW�W����[��&�qd�C1�ю����'�2a���hFų�-hT�pM�U�%�jCn`J�o�s1KI`i�M*z�!��f�,�X��aƓ��.	qj�Mv��:u�qt�>+��Wv��p�T08hX�8��8�l��2�5��w���XgG�fw��+RK�V���i~U_z�����S1��:����}Y����у[���ʍZ����?$9� �GB2�(�yE��>6�ɖ����(m �u�~E:�0!��[)kk��e�`��E�vq���Y��q�]H s�@楨�� �p�P��b�I`��?{+�5K�5Z<.�Rp7p����呢�z�F`�I��?j��7Ҏ�6q��j����FG����oD7-��_�-��w�e���Ҍ�r�������	�� �rL���,h��/%𿕋e�?p����5�Iʾ�ǹ�p0U�=�FiP�W�*_����7 _D:@r3��$,��k���u�}����^m'}z]�r'��B��|P��A��,sX����5�]&�%��Kk�8F�eF�i@W��K�4_�Y(�QVK�������:Y`����+�T����Ƃ	���@F��i���!�5�������@C��:k�-���ؖ6�=�u�Q[��/�}1�l����hmD?�,3�����j�9�ՇEgӕ���ɍ1߼�����V�:&
�����3O��$�D�j֤
�6�k�Ly���3XL�(�FJCd�8�š>��E�6K��I_= ��I`�Eb�^fCЧ@Ǚ��|my$/�ܑ��vN���Mm���6'UE{e���Z��kW���M���j�b��=p!��'���].�"�a�ޅ�%�B��-��y���ۛ#��+ �W�l�|����o�#��(taG1��
�Sq6�//`zR'��'��6��%�D���ɑ���L�t!O�+��U�Q������e�8���3~���5"�z;g�G�?���0^��������k�<�[�	ȑS	��C"�����~����r�`��
z���{�f�&�9���o�y[D���$4%�ͽH�Sv=����f���� ��7�3���>��$��4�x��.m�4�P{�O5[�$eQN��*���S��Hj|]�LT��Zf�=]ׁ o)@�K�dމgJ��Q�p[�2c��xV��QK���O�6�W#��q ����%� �}zc��1/�F��ǉr���蓢11��j X��M:5�3� MVW�[�L�dd�W������T��8&	:(���1 �n�Ft�"1x��D(�{���B��W?�W��V�#�K6������4�řhd|�p���߯��z�ZF�?<���G�O�ѓ7b�܎T[^Vy��Eo�}ԚF���b�p=���O�'�&�E����_!CG q[��ַ�o^-�M	ߔ?�BE.KV����)����^�����^�x�^1���O#�L��uCi��BE���%�j���U9Ш6����>{��@ɹ*ݰ�5$ (>������,�PY�w�÷1H�\/x�<ݧ�[�n�{faԫ��8�T�U	���'�)p��`ԗA��ˑ��� 9��(fc�)��}�J5��A�mM$��o�H[�u������7�q�s��ѷ�Wa(���N9�%�<P�f.��7sz=A�r�x��!��7���(���?�..<�Wُ^і_������'w��o�XP��[1Q���JQ�3�+Qg:A�tC��B�5�ھ��*�
��X��fi�[ǐ̫8��M���و��[��Rlh%(WB����Ǘ���v���w-�w��8�w�X!��ie�Q�$���&1��9I�"�\X	�AG���\�c�u�no@�dq�m�s+%��FK�_� �.���ޖ�=��b����o��G�\� ��pL��L#Y`ѫ2�2�G@2跷	G)6��@cŝV:X$�Ʉ�#�^^P�@�5�%d�Ӛ�r3��&X\�f?U��,�}�5�jzmAﬢ��Z�qʦ�Y�h֢��v}M!>0�7���E���lo�����SƄJ�2Ѣ˳�Q
v��]�LT~e�ɱ��PK��'�e��hcˑ���.��X�xm����e����Wo%�sZ��A�����_5�~���C��ܳ�����N8X����S|��w��K�+�<K�}bb���s&i{����e5H�*���{o���C�$]�6��7_i(GO;�4���9����S��R�EͶ*(���{pr��K�t��[Ϻ���:�{����1�j��*f��G�7�sa$�Q�z*�Q�2��'��v��H�� �����\�h�Nd��]L���%�l'�~��N�p����H��/y�k%(��PbP�������u��亘�Q�U�R�4:	�%���gt�!@��
�Y�{Cm�%�h���~q��Z"ׁ0����
�BH��Q�z��lεeE6�B��We��e~Bp��0<�ρ�~j�-4y��p&m_/c�y����>M �m�"me�*�ͦ%f�)[\�hc(�$8ZtR�P�͉��.��#-B��t!�S|^�+υbi�����]A]8j��C��Iy��O����ᎈ�Ѧ�AJb�.�I]�Q����h��Y�mBu��R���p���#I��Ƽ݄X�D�����E����7O�
��Ԓ������^��s�`��GFr�)��d��!��9����a!KX����B�fy�FF�=U���:��b6��]f���t������ZH-s �QOw�6i���/S?o�lÉ���A��j����H$�z("P�k�Ũ%��\i������A�y?%`	'��>Kۨ�#Ԇg>!����a�-����dp+�W��?��E�JviP[Ý��\���q�Pi������u�Ԇ.�m|�}�0�>����t(rG�1(8-��'u��t�p3'��nym�sAQZ�%�M?�� -FvpM���>�]�!
tαm7��R��ݺ�s�(,-/;ՠJ���lm})�3���LS�94�&�
����@�aP&ƕ\�	��W~�������d���&�&����mQQh[� R�c��Mt��
��C=p���<anJ!�H�v+�(Z/��DD��e�{	K�@�%��=!�Y$`��W��tl|Qh���c>$����0���1�vލכCs��ʮ��ݐ��2�5z�^j[=#M����Z�sJT9��;;Ϋ�6�.WQ�Ͳ�(f�e.���޼���"�֐�a-覃�>f���l/+ʷ���֮�r����N;�����i�e4�]��S��'}��du���ﴶ�g�����<y-��՟�ee�	�����}k��j�窶��	��?���i���̞�w��;��pC�I��2��#A��.	B#8�Z(��	��E�N��';�u�9\�}��s��S��n����ʞ�SVn�(c�:�p��,7&|E�F���躚�Ԅ���LAb>����/j�F�y�:�F�27�����g̤8�q,efR�v�G�y��	�c>-��� �Z��>h/�r�~��H����J�p������B�'�k�������/�����Ck?�I�����O�]`�6� @j�����$
��S[E���L��t�I+���P�ŧ��`3IϿ�U;�U/R�-�5��-�eN݀~}t�}��[�%A����4Cٳ���?�au��9��4�о1��>og���jmȱ��'��=�a�4��md���*�{@��S�c������P�(t]�Xfdǎ�Wp%l�@��vʬ����cz�T���J�*<�"��:���c��?7����͙eVO���ѝ�n;x�%�ɜ�X1J������%c��ῳp=�x{*���,qi�����`��Z�aG���WTf�]��⾫���VL�lk�fZ�I)R��J�Y��Pd/ϸ��5Xv����Ӵ���v�C+��9��0x;8��	F�/ck�
o��>����O�2�q,�J�#q�= ��ϘiV�KzX����{P�>���\d����_�֍�	��2w��K�gh+�b�j�5�Tכ��K�J���-�R';y�6��X'����FbW�'aL�w���t��y:�0�g����_@��O��o(����\��@��"�Cu3����s3]���ٺ��,n$�M�:�L����^�$p����z>���ԍ13�&�(� '�����F2I{��k�_+�%T5̄�x��*rI�n�.��5�eyt��:@W=�ݱp�2h^��1��;�Pߡ�� k�C����2��lpa�2�@��<C` �m�xn.�������+�� �q���&\FO�%s�b��SF~��`�����:�k�?3b�pJcDY�c�su���Q�Ѡt{F��Q.�A��ӓ��Ͳ	��ݧ9��/E��������>�L�VvCž\оd�%&ߜ�ߟ��K@�j���3��$�h8Sj�d���2d�����U��u��c�}`�&�_/�̼��kZ",��g�[�FJx�Ђ20�?����&.�	�Oʌ!d�U2�bq�F��_���U�D(�Z7�6pDx�=������>�0r_�4؇҉��х�Kރ�lh�$pԆ�ieor��E�}��U��V�n�ߝցA�+j��:�� w��TeJ.�CqAD�����D(�����k:ӝ|~�>�⍫�6c#�� ��懌xz���T>:t�����Z�W�z_�Z��EW@��G�.��b���n��=�(�^߽�n뜔����g\+{��y	�YO���l�A���ʒC���.鼧�D0)ޘ���x_��F���-��������'�cX�,`��8F�/�HQ	�!����Ĉ������b�,�.HEe�k��%�� `�L���г�a9yS:����3����yoI�g���=��tmb^&Lژ7h����
F�-+c��5	�!���,<7��:F�"Ц�D�Pn�W���r����l��e�;{GwK��(|ePG�QI�]�L�Z��v��P�� �1|#|�'�P�o�WY��.k9�}#m<��dM�p�P>iS�C��W]�'!O�c�] �5��J��˟:�;.щB1]������#�3s�����o���s.K;������	����8%Z�B���/򆜞��fO�6��Yq�F�������ݍjfȜ��k�vl����]7�$r.+k�Gґf����VR���5$�v��'8tr�	v+(އ�>��re�1�X0���a�'s�l�x�/�kO��Q��?� >o��47X'i�	���hUe(��r,@ھ��3�J��$w<�\Eq�y~o�jo�9�\�ܦC��J	A>Xn�E��UA4Ⳋ�y��z��,qJ��Zx�T���zv����v$������rW���*�b;*zy�7?�����FKo+��HG�%Ip�\��h�AW���é|ؾ}��֍j���%B��a�
eS�H��e��H�֮�l�Ǉ�h؍65^�G�X������q�k ���DNĞ�b/�x��������Շ<^��wrdzZѱ�������kNB1�5�#�Ӹ�u��������+Z.��ΕUt�̭��l��N���,DH�yV�aP���-C,y��W'/��Hf�(e�c=�A�V���ΰ�"b��ފo�Q���JN罖�6Xd�8g��wܳ�(�QgҞ����(p��+�,��*���?��Q��\�9'��"����&��F�A��͖���~�%㰺%��?��Tt���1�T���XR���x��������eî=׼�����1K���N@�+�ǹ�fh��tx��Hׂ�}�JUrI5�TR�z ڢ��}���M�����;_��*�
�Nut������>>�Ta��Ijw�&������8�4��"�ϐQ�0I�5&{s�2!�*�	�ׁ��밺�ű�>ќ�A͒���_) �b���4�7����*	I6���Yy8k��oŽМS�VfK����sH�̯���c��-$/N�]It�H�.ɧ���b��A���@�
~�)&éM���9 �@���&�D?�9�>CL�)�3	���C�D�rC�#�����&�ȟy�2���y����u�
 n>�["#9ځM@�[�A��j�,G��4��%�]����t)�!�,l�'x�EA�w���7��;h���F)�&-VCP������s�)M� =9�f�.�`��'�4N�r�1�Ө`I��7P�b������v�Vu@'���a���kazU������}y��'R~ =����ee��_.�M��E�K�k��0�ۑZy�W�\Ț2^��ʝ�x���e'��͒�4���?��r�̜5����mh�S���7n�$��M˼-d6�B_�@I�E8���i�E?�������Eպ����*,/w�*o�Z�~r���1��1KI�bDM,������bx�L|D�U�����dioN�=��+F��q)e�o�\�F.�W���a���=no��(MKh�������l�i��"��r&�K��GY=��lf��}v��A��b��3�M4��0�*y�H��<ט����� ���y�0+���:>'�`J��i#@�{�U�����P�]�6�������Q1���͚&%VΨk�#\¡Q>Dm=�J���.MW��k��Qڄ��ʐ�Ԁɱ�Pꀽ�h���J nS=k�fݵ �}�E'J�!�!���ޭ3]�y��q5DK��_{:�a�����t-1h{%��:
��;��I�驑bs2�RyTXM������Qo,�P�U����P��}��6����5X������(�nІ������z96X�)��\{��ygW�k	;/pڭX܏6b(��N8xӊ�c�Y���/`M�?�>���R�"\�*k����K���+]�tS5&B�0蜻�5���g�@�������iPS�D����}jo`� �1�8��xT�?��ޗ�)K�|��N>[�NaQ����b��.��wM�ݘV�>j���d���,���^��[�n��ߘH��|7'��mRL��ۂz��[��p[��u�r�w���RLY�k�65��hX��9g��$�.�	Έɏ�v^�1�/5M�<�n��&Q�s�����FN���Te���6�J3���8<!�-�cʽ�:��~�S�cF��K��w��Gd������9���vMG�<C�]��ݖy@[�y�(G�WF]}��C�z<;�8�ݪt��Aȁ�/c3�d�,�;��/���ڋ�M�1�l/��ru9��*�w�/��'�i��+l�W�ji8K�H)?Qއ�T����D����KI����wݾ����Н�.�%f"�lC�7k�w�" !W
�]Sz�����Gg�.����(Ob���8�;�H`LE�<��4��:<��@>Ax��&0���1�g���y�r��x?�_e����?�̬�3���3P��D�:'�wDǗ���9jQ��
��T(7��#,%��y�R��*&�����!Wa�'E��\�}���ؑ�ZS���ճ8٤�N�I�ѬuЃs�d���YFH�xWrw�A���W�H�p�M��LDp9�OZtC!���QF��N�;����.^�&�����=:�6�#F�k�3����VO�G���<׏���� Ӽ��Dܟ��F�Bp6��(���'=g9$�c���4�A7��@�4~�g��AT�#o�8� 3EY��3V��#8��yHV�H,��#�ثׇJF��F�!��i�T�d8��%��߽y��H4�*D��[��Ȁ�b4�NGEE��E������n)v�d�:<,?ϼ�� ���|�.��
�kN������%�w�*�Qq��w���F�����o0���:���kE���c����w#����S�e@��,�*Ĥ�禌����ꙶ?K�����є"���v�XGaC<��-�M�Y���`:"�'�ě,�����	v��䨚�����TiS�6g_�1��I�O��0����#*��E�R��S��r��!��WMQ0�n�!�hj��?[�m脔��
K|�nԧ �����y�gt
Y7iƥ�˭	'���(����(���{C�FFk��;?�F�0s\�u����O$�<��Y3X�[@���2�K�=��Cb��D-J~�Ixa|=#���(��.������~����Y�����b5\H|��?lzXu\ C ����4����as�m8-o�	L�a��?���w��I�9D�MK��ҿY"��=�{#�k(�K1�@m�b��*fu?@�B�l�GiKR���	iu%k���,�&�Sh2�Yj�*����F`"����gF6�?l�cA?�vX4�$e2b�ت$[���"*��L�Aw�o�\�w�?G[V�R��$I�ǆFKrh��K�h�BT�Mi��	��;����B�`D�mX�-s�B����8���o�^a�-���|�<+T���ZDdf����=����5����˜/󧇞F����1�\���*VuЄ��:,��tC)�D��e˕��L�t_���9��)�~��4�����l�XF'���rqP�UVٟ��r{��>���Ek$��\%�]j�� 5-��irӵ�?��ǁz ����b�~9|�!� �D3B��(U�2�2[ώq��6�3� ��@�i��z��(1��9�8�[�E������d|Ϙl�mו��P�<��2���ҿ�r�s?�cL��X��}/��N��p#;-��V�I�=;�,���XrK��m V~5K\%�S8�3Vq�9�����j��譏��j7ͧ���k>Su�qr!������?}���^���z�u����0�A2�vi�K~pý��*���X��CnN�3T�aʣ�Z��:B���ͧ�QW��t
�_+�����a��8�+Ɯ�|@&�x��&=0�͍�CPI��w���L�Y��\|�6tj��c�HLnG�'_��t�WfW�_;k���s'U�ϯ�tkN�� �?è�/��>`���7��:<c����޶D��{Q���R��ՉK�G���� ���`��L��'��Ԑ;�):���=�>���J���x΂�ч��8E��h6ѱ��M��������P�6dݢ�P/�������?��~����E�&��X��h��X߭9K���Z��pu ���m�/��[kўķ��Hu�҈#����~vCR/�:s�M��)�}ٶ/_�3e����i߶f���g���4��)z�F���I�k-��k��p~o��+M$l$��\�ől1�^U�=S"�o��[_��BnT'��8T�O��o�ўo�K�e�"��.�N�g&(��������'��q��XKӧ`���DRK��Gg7��.2���MKn��@$E ��	��/���Eq_��y�:w�@8t���ո���+��/i�n��P�����Zۋ��}��� f7��[b&�g�畣��T({�ݷȹW)bAD�7�(LꁾL���Q+��ǰ\[�d<}#3�p�6Ŝ}�~s�������