-- (C) 2001-2016 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
MzPnmGWHH8UfUjVqPxr8Y2Epuj/asSur9WqVprKxrHG9Cu7zBhNacd5BFwgJgntTr8AwVFtJUeOp
LyUu8jNwdlrEvficWkIHGMhvpU69YErnvwUtgR1mrN2Di15uK9rHzl92BE70AnFi7C0sWIB/T7pc
FweYd5YHI5fv6NZk37i94GKWNN5uSOPxdaVM4ynZGZGMN8decSNMV0EPh4AYGRV6KrbprNoa7GhD
ICq2J266lVoYzbo7jXqkRMxbhJId8PdENKTCBgVuPhlcyciA1w1DtD+3WOZe8vr6XXBGbNrFVSD6
de/kTXcNo10Jjqkx64JiTJngijFaS+yekvsekw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 6784)
`protect data_block
GatwyZ7hjp51VwU+Q2aYlrtpAE+OtpIVuC2xVxO6KjROvC+0oNDbaLhgBkU0bxYVcKeAit1KF9YX
jZwPOdaSC+n7ByIMh6G3kGHa/BV4GFqQtDyywGgvs14viHDnMqwmM5Pku1p4wynZ283g7fF/MNTl
4W1hy+mVkeHbAaUSkJlPLOmLbdL7TDIqac/RCcYIJ3Y4yfwqGiiSKaDX9OkuHTtRNm9+2whqiRwV
1R+EcAPTGWNxChFb9+juZ3yuJqUXd64NsYZydvbncshqgAorYHGwd3QE6LOwwyGFxvBnBjrF/+Ds
obgwza9JpMdu7P/6Pn4yacLfu6rLOFga1ffjcEJDeGIlL5aIIhjd2Ku3mx5TjUWoozyGgn3s/0sm
lxEHV1s62kkNabjrcnfn5O4pWp4Z1JRbt3v9rYn0pP/8jmSz0pvVVifPEskOaUtI8O1IYzK8yhP1
70f6LMVYTI/sFa8K1JiGEMXbqeEUvxKspUUi+xns6EXsJPObEonm3Epiw0SJ3KfqNJbIXD0Z6sdE
KQDCrcnOmnW5jpeIk+Xxu2Z7/D7wYsNcZzqDc8yrMripyyUD9/yANA2FD/7QnXgkUf+S0+wJwK5f
iIsF9xIURP0QM5vFyv8iM87vJWCEBQ2k45XaOzNc9q7+7K9QcSbELkbs+WTOkYQOsIq10Z+AEWis
Karw/WWxtxlcju1NvWp4qhlc7WYUF2ZdRQmw3Igh8RSeFTOgONg3sMbMR4ztxqucKSrAaMTMAK5T
NIsElsAQCgCGsCa9UutMRf78ZEZ7ptTWvk/y044Pok/xCQZpw5K3dwXHdgoJqjNs4z18nnm11aOz
lTeocz5sVa97Oa0BgCMhkn4GV7nH3iIsvy6z2xHSbuie5ktjzs7f0CMbC6SWObh1kbrKsnoL9Flt
iwkZ8i1veuhxNBhlKtzLpzwT7e/6P02J1zloo3c/XKLfpm+9EwBR+GHP4p/6r3TdostiRVAgnRZV
Mo0W6hGptyoGoXIGTp4P/Lt1+BvUwUoSVRyutwA+WIwFII8EemLSCHeS6gMEK6+U8RqsDaK8zm78
7pyhHTnbnWaHgRLYD1BawlzIouZkQM/jGdUwATLtTPX14rncmMI8wkBFR6v8HWg4rGInx7LWiaXg
qEkQIa+9AwTsbrEvF1zAWwdJWyHL1wFleC50i2ypGR74ByiPGfrRP9PxHfBW6Rjbk55I8jG50bjM
TK3Pm/vEczJU7z1HN3JSQ3/3droa4ddOUc79ZEAUUqKd75xT7qFafZxd4so8hslsBweNt6F3Fbvi
1BDPP8ZbGmRNRg556lVwSMigJNzvgaVO7YWxOYut4badHN+R56d4j4jg3NtTjACsl6j/WCT8UXtE
ZGD/6gZJzoRAg5MD0/26L3Ueoxx8vD0T2mhVsZJurv7wjWKMElwHfpvM1oBrfPcsWY2WBqV9m5tT
gk82IX05G1XGY5wNymwckxCOr6OtC5YMsHfluoRQs001c11/FhRiIbRyZ7RQ3bkyr2cpXy8ybqqX
a8vRLyK1opd8++C0CqSS9VxxqzmDtndmcnZUcSjVkLomD61wi0bGE1uVAONfCaiVFoT8rygS26hx
B5y1qZHdVgAbMvWgcKHjwDQpdIDBLaVXTyYau1vYynCoce2tDYQ6G4yRbkjOf/81NuMijyU9rL0G
8pVoiojxrHG9Z2ExzrMUUVhdhBBonFMHwdWZXsvX+jCVhv98aJKu+EKcDjLJQ5jD19ciQFDo/fex
U717oDk7/yZja4zvSoxyNrGgxv6RWURB0p+eLEoDG1iShJaVXz2WUT5/JJUGOCovWPaBXClN+Lfb
d2TMRyXvU7IUcCW0Kx75x5MxPLN23Mn+cou8Jqge1eHeSLKDfe5q4BRMknAxwivtvX8Xu0N8fcXf
5yab0LYnEIwisyLPeTt4R2Hh7nFh/9kfRhcZgW+GU6Nw+sqnaApn12JF89A3v6p299WPiN6PikjU
/QpfHy7xrrBtyuewU4M2v9w4spOxyNs2DklfMyUu+weVjci2yMGsTL5fvSg5KZvAympIgjIvlQOf
wEC3eOndxb7xZBIDXdLVWTwNLAfYXjkk58HZTp77tnUE0RrEIwQR0WdOtxhqxgjQyayC5+UKAjGH
8rLAdXNXj6g0/57p8oT+mAKj+Y45CiPNwXossIFP5bScbACrKrg8m9oQKa3DVssbLYWI5MJmJATc
c6FavTL2dWP5j2j8V4yvtSWMY544lUFc4PjK0gO5FfKJepY/agHX2ekwriSivnI2Eiu22ofUd8n3
4ptaWjFgzigs+ROo+fa3nOO/UbEAaP1/XP7xxvh0lKnAMmd3LsOFA0najt8j+WM+hPKXdp67KTvI
QVo1nIIQNqH5FYaxl6KfvE8IdRPCZuQs2774vTR9GE+eUOiDEvyfXtS3DB5pWYOnCE6dFSQkO2Ws
qD0hMqhLyEMdS5zxLsSKMzPDHWhU5jXdKhg0d5KTkUEk3Wd2jOHrNU2G9g6Eao5iMl/AIHtNturc
YBnBoM4PftqtiKvKUlxEy5gxHEQMySJLP+m47c137Oe5i1vc71KG209YLIivaITsbTtkU+FvkBz0
0b5Q7jAFMUs3PGYcaEO3N+es02n2MTxVaFrldeaSd6oTJmcwH5elE25OR9rHQUm4yt7Ie+mrG6S0
UxBqI5a5zMpuyk6ZQ1lgYS6HNFnIIafDWFLdl0rH09pN1az4I3EOAvzW5inpVhQ2uw6MoiT/fbKN
baHX3diW/1TQ8Mtfy5nQW8C6nl0Q6uhRxspr5wvQQxOyBE65C0n8QmYVoJSKkzdpVNQRvg1p1++u
CK70NAbVOImAwsrw30khpzvxKqWeUJ4ZZerDAsooV5JoR/jeWZdCT+oqW++mK6IsySrsJTFuf8e2
KRXkwPd83lG1KyQOtNIBfPV9pusIEKlxkLyzvb9ZBJORZ77FzU1LlrLyHaA5G/vVRNf+xW3epoYp
S8xkIuswslnILz1MzDN2R9kySTqzwzkbUh6xG1CGe7SYSsL1PPFV5RAygcvHduFxhgCG2l/fXqAY
kmggiMRSFd1I8zzVTX5vb5pMqgI62AO9XBOa7UbAHeL//dSfDR45atmzlY+YF9hiXmU9HFFaWp1j
rN8ymmc4K1EZBCfkRP39QR5WNKRem1YEeuoTLBKR8hWUpm7qmC8mSyEG6V6oqeOztn0FW3oKDQLK
Mbe+05OqeLPNmpY1OG3VX8dKNjqGBjerROcxVjocIoi8gffyIssAmFGXOfJk9/lWsl/abTWNaWp2
A+j+ctWVZtastrlk+CAgIOyIaR0nDbegzXY7NcdFDR4k7zyfS2W45bSZx4hsQnskkebDjvUbkJTM
Te6wT7J/9HT1hvTgw/ZeK+WCT1BPKnasTCaOWCV+QTvhwijIJFfQDDHVdJaf2MK4QyolIY289qgd
NtiYSV2z7g0EeiIfZ/jVYNiP0odai2HS7oz6wdu1zeTxG2PxxZYZVqAqJ1m8qK7UJK9gXTTXK4zZ
pJCZqiLkgUOQgOcA+cKRoREY7/+nt6Dxr4ld6ADkuo8yh1/riv9/OgVPh+22XTef6OSbzZKvHzXn
EEI0KUPCNaJTlYDWyFipNAiG3Z3axgCJIrmLVZCbg+iUlOZZKIDs16lEsKqAgz1aJpCfIYpd4YPp
PBhKszn0myNi26FrRDQNJUPCfLe89yVEaTSl62ThDSRHDpyXkieOwzxapx2zt27wGIw9XxEOn6e4
lnPmc8uLvMv9G2kNJ2Tlz8ISjXT3gzQcIMrznXqj4H4BoTC+quCzcTtm6Q8u44uExrrhavhRrfth
6yWUEkM5irIM37wwnPjacnWxsq5LPtryiUWptCqPLHW6AXtD7+zeZstacfp9XO9piEYnGn+H9hAY
UufFDi60ncICGRDNCrVAZ3zjRFPmLQAYnNX5dZG/eozwE2QJsB/hgKAFmF5Ie9tBjl5Yize3qv27
i1oQgOLU5M8+3XwGl8QXVgOTMYPESuwtQNzu6isr9D9+liloAKZ90O07iMPNP8Q+JVi/hhXydZEs
9gwI2laf6Jwlt2nyrO2g+acJusyvmyb86mn5fjzxO1GBSWUzonyDDRx+ZirRfyP1nrPuzuud1tgd
55CbEAoGG2RSyecZLa1k4B7ojVT69HsFB1nPQnljaf65m0CeRjDBl3y6z+x8iNyB8zjrLF4Pbbpp
Hbx0upx1CfGDi69koyDLf1LGf2DsLjqWkSiWi4mLzCGwFp0SjhrzCmk00gOFL68qr4fGYeF6/ik6
cg2uEZu3qR9FRdVFeT41n8981qV8ecAJn+NHYaWzHs55S+WtqRhYdaNZlQChGlq0yHcYASUViJKU
EC8Inp8Ef/vw6CLfSaCsGhPfgtRUL1oEzgUhnqcvnXYFJ2sO29NLz6eTrXTAVel3m47YoSJZHHeJ
/qlKPiXrBdSFq179NbkgD6de6Lho+Xk30wwX+DM8XsN87S99CERro319gtkGoE2YOb7BgNb7JGEc
SyE+HvBcORyivw4wwY5gNs+sSNC+W6gVYQBSiv9VRP43qqXbmOF8GTaxXuuDENPx8q1xZDsSMORH
Gtrj8cN5Ufz0mbqMU4A+t0QgPiRWzwGGo+uP8I1yIWfT12Bufi63ToXNnNU8ZEFwWh96T7ypehra
U8niTl2f4gV9G3/eSwDF6l0/P1oGz2EDcJJcdInBDIHjMAJSZwpQuMRQwnKzPz6ke1cToNAcM1FH
d7skx0sHdRux7MHbuM/E9dLAWRMM77Bi4kKhP0IdVyUdoXE7w0iWy89l/AGM9bjwxSfqTSC/mc3m
NQpkgHkafopwqiRj/VEwDakV1Q+fsXGUaw+JCGcEr650J2JLjksySmSdlrOfk6xF0Ti3Ss2g8j7g
NJOKpDLE4P3ytIVjHSWQWgCtrwSAJ3iCEEymIToXewC6eHsR9Nph4inAQCUEEbSYF3AcZxFkRuq4
uFZW0A3FaFFFadXvoDcgw90+u9Nt/nUDpFBlC2ZsmnaWljO/okKK5XwPiP8bHX8jCq8b62qQm2oQ
u3NmDfp3MaBmR2bFyw8EWlzNYiXBfte46MlIdJEvG7OktSbaIyK9hhS2IGpBFuPFjssM+1ynZJLf
4e9/ATlD+okASd6lLHiJQdM+0k7STXLtWFjBjJhiNHDDxFBV17nsKs5TCsD74iE8jGBMWMo2Q5F8
EJa2KH5MNcHsM3q0kyH2evuDyZ943nSVYD8uRVzw9gsNcHTeRAZEWp/d2JiVf4DaYP4gku5yYMZ2
k1FkMwPD8zNv8kxCAcQrOyGsiRHlkaSqGtrjLTjwUrIFW0WvfOC5IF0RSDbFpUWa/625PY5RWjas
kkP3r4D9fn+DXT+ZmPnYLEWfHyvP5dTqDbbdqb0REltzIAp6IQ7vn8h0wT4h40n8YeyTODmGH3z9
Pub5baFtivATt7ZExCCLbqcqXii+wkkPUXX8zFqkNA8Cs37tDjkcT/k4ZP0f00D9MiGo/rWGQOJu
CIwGVwqoYx8qi4Vl+BPljJ38zkffCvu0w4E8lzkwdtQzuFBZRBhL+X+i1JBrcLrNnclLKVS8+zBJ
1oAfxZq4dEBcBSkoySLfXoUJRkVtWSiIpo6TWp41EcAVb6XnfYz7iSH/ogKz2B8DmG9j9Kf5GAtf
VS550HIeSCMbdCehNCRwTRoq35y52ahnSA0Z6SFZ6pAqzEvwCgI6qHa281rC2Gmh4NFKXk6qWiki
B8TtYfsAjQTRXeVi61CoV76ikpt2nGjw8uAx972l33rXUqjd2k9NJ79OQlOWFSQTg+1vQbLRdveb
4raZHBMlO34tOvceP51nNvtYgyh70xCQGPleowPwWS6+JVUycSIXxGBLZVQSzmykkcM1ntRgGuDB
wVc6dXfhOMlkU9W0TPQIwXSCvXkdpL5f3hK2cTBMDWop18uBfaUSAxbDj+OUXRoVYcOsd9oy+KfY
Jhs7PHfI1vSo32Mw6wV2Bg00Ny6J9jRxZbbKGxEAlqmcunyO/Ggvjpb574/S99uO1zUe2RG196tQ
Z0uzqeakORDtQgdIDtYCCrwgvxKCNtczc09Qa1QKW/KI2cTeO1porZhMBzCe1nXOid4/lnOPtycJ
UvJuiB3BPd+1vEGAfRInQRd85xXQ2tEmOup1y9lSKX7Nu3y34ryp1gC6LLCTtBNws3ktj+crH7xK
BltPNnObdSNJOLBlrZhcqzASgP2Zz+dv/AHG7PmatnZwEJasnZy6v7SUItNLgDncp11wGaVkdgdf
njqEUkpGODEvHAFAFx7AMDgeQ6fjZhNSNGGmdRenoUV9Lv6QEzDAmllODJqyY483u9K3BWpgzpLL
I0vRcE8FDaUPhb4iU2YeAySrln9HM6H7WvWn3h4ZI4E7/ny2Zx0wBTyFmbcwqz1hv2hsOawNx2Ek
UV+US8q5WbWTnjKxm4l5svCNV1kwrMq8SB9e6ruT42brO9KcPHzIjl/TtT4i8bmIxsL38KeRFIU0
+DDKdKwXK+MaKZWkplqlXNUoP8Rjk2MuYcPjo9sDaPh1u14G+gUccy7GZ1L0WwQswREScVLpib6m
+NeQyIDqnOC/69Npx3ZFu3hVUhpxfnl9bpyBhat+eUd6VkdxPs9CV1Av+younEYwmhD00mUawPbD
2IA/L/HyjvbOIgGcV0tcwGWrTRESsJYGk7QmO5jImUXf/9TMtImSJ5p5NcyaN/1MZdX0FVqs/njT
OvvAd7yAIXobtDpBbL7ywxk/u+0Ya95Tn5GHC9YfgB7QFLBxcCSRmJZUqOuIAn7/szTSEDzYvNjT
aaknsNjnn1JBncehmgwS8AP1u3z588gfxHkH2CE1Jt9jprFIu4+7IfI1q0WUhWK5pDR/kddwaGkM
tl5INkZG7yDEA+DaqhFMi8LZiUQguOChdFvfx6dIXIQvSnx+0Z2GqoK7w05CQdTBkWgtVfnollPb
Jl8p5uTFR2srDRxtt/Hgaa81FSsIoIxvfD3rZQThTDUSpHuPkUrpzcHRz21iJ/3YPquzjYOg7naV
ZodHsiJXm9Uwx4BRFMYheMkktgjf7ddXgjisIJF2Ro9xNWfw9UWC1JL6YUl3aTG300MvcN3EjTEY
wgiK3oY92h6foNPR660cc4bYqYOke65FIlk3+pXZzLeQ+HkBT9hidM40YEe07ySTQ4p8IyHGAzF+
CxKUFV68WIPTGSK1EhTUae6YE4a8Q9/Hy50TGOVi2sx8M6+TR9QqUC41h5qiHn0Y8uy5uvCYDSDF
Q3iE4wAk/MLnoXJFVIj9iFpRnYYKqoRCCPNu8NQvvpm/X62kQ3JEacUR7tMCJlKDyJevUFtYcMWG
6DCchT2y3r9pN3jhRMycsRhmYU3IGExYREDRsUVgBrnrArwyKshKz5LeNrZxwD2o2c921WNi4iNj
AW3Mb1oq87/oWw9ZOXVelDqI34XYGeFKmJo3u/QaNXGw2NoZkxAryVcdhQDpQyXiiJSPrw5giPgB
qJ9/1CcAZSMM8w4KFLmvVaeMrgVwjFs+WIchC7lBN/OfBqnBhdGFj6aKeuNCZg0d4B6TJ5ro7nB/
1SQZbQ2N4HzegrTrNWbm7AphlbWAJpVy7nN+4fqmIpwar+SoPDZ1l7gnMxMP3GhMG2u/K2aLHbDc
IIOhjfSLa5ospiHl54Z08lu5cjg+m8IhMQ15VbB8WIeNCrEpMrcsKrZgr8l8Sq8fNspcEZ7Fuvyk
KnYrm+nYvkjsRtYHRuY24+2FpT9pPQ5gHtT5vBOBUb0CgGvfYR0qA3qoQSBdIrFfytBU9fscyGzV
RE57ndCeJv7JjLfweI53C6cYeOodASqvI0/Llr8rVHuzUtNfxST3PCTHR/lsS7x+Fp22iueV880d
VEPrUSQbduNq0O/kb8B/OPDu+2QzAFxjj5FniotE86oNBdC2+KJqc2JMcTcWP56xQmW5W7Lvshth
wxLQdoEwHxbaWi0WR44SixysGKylj2e/JnQDEtzwtkNp+88r3Ag2n7X+IN5SOgyJ89bYTemQYWac
qKd9rayIFlmbEtR+yQ3d6s06dnxImSN4tWZlyzBJsP9IrD1ttoiERp3Mmc3uL40gb4TRkUTZYNmY
w8kXK9JAm2XzyufHFTVFUYh8PAXqCVymu6bEYP6EC3CAijTRSNXymO8syiNNAPZ4qvkmEVnwAvwU
dZ2bDSy7OwzFquYooim7LYhHj5HRjy3J7+aYj5dKn6qc3Q+7t77M/NoivBAybMEDJxdJ6A9C6c+6
wHMzcmZ+1nBRB4HvDcA8QRHtLtUEQ7hFJIYnlZL72DQ4NunJkNi8cZjAD60Qbb5UzvnW/LZtAUc7
/5lQleH/rSiqGl4H0RGs7Ild3IgScf5IboT/CuhCjhjKEm4zEVDK/nqb1puaXDwNUpjXilcXAowp
+TLr9A0pSyi5S71FgAv64EtplL2vu3EkVGXdElnX3zAYkTQREU54a5rVWpAyzqbILIr3BWOlHmjL
yB9HpT9EMyuUIK8tR7cVWY8ASa5sVFC8oDUpSREyZznXhOHjdoeAMfSdXHMRcGhyPG0TgC9yI3Ww
oC0mhfXvsLcvxUOj+qIXNp2Jg0he06NT3XgFNpSV6BLVCXXdecvxw9qQxM3II+xHTfJ5SDT58+o6
IlmPTxZGoD+3rAMfXeXS1pEJI2gmJ9pom7eoVSVS4an4IKWyI7nVhBMqu3mBzpDoa0G6EbvFruCB
sh1YC8zQYiLqGA2YWngmjdWUJnhJV6Z3x9MwCQIWQfpYWRNo/A+oVg0kEoHDqi1Qb84GBeztOpaw
7/3+yT0aArGKNSYQoQ5/mAShH+D3WHnMcPQYb/LAHyB6vZyKdU8uWYliz5LZDUAWi35wNtkXdv8e
6mOi6HORhZ1NZhKa+9EslY6J65vXUQiAe4zHLwwZzmbbqHwEF20fP6HOskTGI5AHu+c2wPf4RTNQ
k4OeISkgy/KLvTJ4QAb9vlf5Q/43f4ArSkQ4zZMtl8US6wNdhizD8Q9GzVPHAeYmHlfQ3kobThc6
KcziTwr7p7Yp6Zdfd+hhwsCbhOd9OBAoUrCaMT3IoP9U77dTjNXE82BqFLUO7PGjUgu0kRFciHXq
PA==
`protect end_protected
