��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��,�y�}�ǰ�=4d�H���`I"��W�`r���T:tB�T4D�m�)�	1��I�t��
��8(�8t>s)ו�."[�漆���]�~�]��;�O(1#5�-� 偙O��QZ��~rL'�x[�i,mׇp���O�I43��4d�,�H�����SN��d���3���r��m���̨T�I;uj2Y� Er�*p�Q$Gm���p�V�`�2^���,hz�<p��l�Bxt�5��s��\yq���#�@W���f:m��T�	,*�񞭋����_��㧋l�	�\�:��uGd��PǷ��N�I��_����Tuv� ���us�(H�~�{2H�:Zor�Q	#%�3ˠ!��iS��95�,?�.���/�F�i{#���Tp5����Ҥ0{%���2vpn���X�����@l����3dc�ק�3	�Ed&3�ZN O���z��s�yxӡt��v*}ԫy nj#��lc��m戭k[��5)�A#�����8�!�]�Z�s�M���t��w�!��'ÒE�rv��Ϝ�c@<U��\tq+��&|�&X1)C�����r�A~��B�&�����s�:n{p��͠R�X⺂L^��R����c���f��J^?��ܣR�O 1�rV���:��T�4���AD����˩�F�w��)Dm�O�b,�a���1$��c��7t[i2>�ޔ0,S���󧇳Ϟ�ᒨ�-��}�!6��Jyv�醊�^_�(�H�(y^����o#����X��3-�k\8�M�T�"`R�DF6ȕ� �,5�;Ҭ C�k���1\������k�t־9�}���� ���QHF��"��t�9 ?��{E_�7��!����]���-�p^8�3 ��TLM��q�"��z�����`%F�zU��K�^�Y;FI�$�*,���!���w~D�A�]�#����u/��eס�yl:TJ�a�ȆJ?fgu��!0m��r^ ����=n�u7�	(�~I�3�'�$����`A-�Ӡr��~�"}[s�����x�0�<�|{�NP��F�t����A�/�j�||>~1r(6#qg�5(����c�i�ؤ��K��d=c֓�98��׭��
I�1�w�eb�E�`Q5�n�Y7�o���Gʣ4b�Cc>1�6�0��S��' ��o8����#Cft�רΥܪz�S漸�b4�QB��|=���j7{LJ�V��u��N�Zk|S�S�=�6�=Y�B`��K&{;�T���svc@u�g�P�{�KY.3���1"�K�\P"�l�N| ��IL�jQ����W�0�ytl��	t
�Te�8���3����Q8�ש����\ޅ�j����Ѹ�}�i���O���$��S�D���a!���W�O�X%������3]��'���4��Phe�cv�ÆP;��0:}�G�w��䬈�>OEת;@n����e"�7���� |"+�I�duG�W�5����G�9��5���XW2�z;(9T_�f��E�+%��gP��)�W��p�>�'ڊo��NO��L��k���������!t�u�%�r����v�	���-���L1�-����'�� ��5 ��<�X�Y4�+ӵ�e���7{=��	BV�7.Y��C���l�1݊��P�/��S���a�Pڞt۱��
�^c%c��6�7=�Y}vC��ߍ��l`~2(�x0o�˱�����Q���l��rI��~�գe�
i�	�E�����ͧ~��%����}�ƨ��jMR��D}�P֡��)��JڵT;+c��qI�Ͷ�E�V��3�����r82K������eC���lD��<�Uޜ#sqؙǑ3B�J|*)6|�����KZF[��<LzZu��z�Fxk�	��lQWvkOrQ�d��d��wf;8l��
s^Y�q.F-�F7!�D(7�yд����I����/>b�v��;G���49�H�`5�U� �w!u��r�n�Q���<B��5��ԑ�`�:l�/Aa�\��,Y@�!�עM�3��?{GSxbH��Vv��X��7G5�� JiʬJ����Nm��V<~TaH������y��w"����<R�v+?��ʩ�3�&����&ڮ���2,��
Ƚ��}�S_5K�Kl��g�0k�����1�����Yk6�Q�40
���!&x��p�~
NL�c6i���IC.��~߰���\\͆�5�=Acu)�"VKQ�`��W m5ꄰ���ִ=�V����������}����BH陓q7�zW�'�����X��R�;)�B
~5����������!�����k��l�TTǲn�gC�<q�:QI��L�Bт;����#V)��Ǌl����3r���W�O.m*N��~���zj R�
��t9�ƱV�%�擿3e(6�E�(��Ar�rݣ,C&�V�\����;�ɢqxaI�xj/�����5�aJ���+�c�t�S��@��6�`I��d�~#���kg�=q�����.