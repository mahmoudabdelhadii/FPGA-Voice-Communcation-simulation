��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����N~@#�k�0!����+��=L���0�ԴZ�2�Mc���ZO�����=�����վ�	"cqw��a��TS[��{=:�����K��-�մ�(��k��N�-� 偙O��QZ��~rL'�x[�i,mׇp���O�I43��4d�,�H�����SN��d���3���r��m���̨T�I;uj2Y� Er�*p�Q$Gm���p�V�`�2^���,hz�<p��l�Bxt�5��s��\yq���#�@W���f:m��T�	,*�񞭋����_��㧋l�	�\�:��uGd��PǷ��N�I��_����Tuv� ���us�(H�~�{2H�:Zor�Q	#%�3ˠ!��iS��95�,?�.���/�F�i{#���Tp5����Ҥ0{%���2vpn���X�����@l����3dc�ק�3	�Ed&3�ZN O���z��s�yxӡt��v*}ԫy nj#��lc��m戭k[��5)�A#�����8�!�]�Z�s�M���t��w�!��'ÒE�rv��Ϝ�c@<U��\tq+��&|�&X1)C�����r�A~��B�&�����s�:n{p��͠R�X⺂L^��R����c���f��J^?��ܣR�O 1�rV���:��T�4���AD����˩�F�w��)Dm�O�b,�a���1$��c��7t[i2>�ޔ0,S���󧇳Ϟ�ᒨ�-��}�!6��Jyv�醊�^_�(�H�(y^����o#����X��3-�k\8�M�T�"`R�DF6ȕ� �,5�;Ҭ C�k���1\������k�t־9�}���� ���QHF��"��t�9 ?��{E_�7��!����](�S��0�q��w�9��=�i]�1�GʦȪc�W�XC�|�$��}q�6����zf(����լml�dz������*�eLD�*�,�m�]ہ6����D�Gw� �g��' A��)�m���b�����L~�B�3A�/15�s�dm�\��rbY�6�g��x��E����Uf��)
^fd���YaŌF�<����^ڍ�-�L�A�hm�Z���JA�&�拏Ӻ�*�=�#��Po��[U�Ƞ���>�-:NM�)��Μ&�^[\c�s�.��i�����+�G'Y�h�8�|��d�j�?v�,�e�Qy6p#��w%�J������q�O�U�>�(zHO�r%�`V<�Q�O�+�Y"��9���1����zlP�
�#�i7`Vq
|F�L�-��x w�lP�)KG�m1�V�Zq�����"������kjk��KxFR)H½s~���n���0Υr�\��F\���(�Cx��:�Z̠i*�TO���an�2��8uꊹ�TLGFz|2P&�F���#��)��"N��@;���sDhʌu��'�GDrsZ?�(�[(D(\�"��.�7��~L(���g��r�=o#7Ϧ+/�~Nk����E�(-!p���z��=���%�'lO�]_���Sɠ�������%���� �x��"K�k߮�!P>� K��^�1�-
&3��t�u���LR1�C�x�c�\��˅2�!y���9�_ܹ^����N���E���C*Ӑ~4���Nb M'F��wBDd�ڠ�1�݃��_�6v���m��W�xؙ����
m�K��1��}9�-�e�� �8�;�B��{}g�l�u�2��B�]:Bh�� �%L�*!Pң{��@B8�T?P�h�-n�+�Co^M(�U�Q�i�g5�
`�W����7�rU7�3W���[r��chr��P�������|ϴ<`P��!� 	F.Ge�Xǝ
���x1�1�24����V/#^�����8��-PAG���c����w�!�Õs�#���q!�Gȷ���0������Nx"ƺ���}m�r~K�\�v95U�mH�t�b_����e��U���N/h4��A�肸��U����s`�4���Z����c�	<{A�ie���k��׬� yf6Z镛0�2��������iˢ���#C��U��0Z�c_]C��Z!���jݚ1�r�g�MJޮ�0�i
�4�³'��9bX6ʢ���-���7ޘ��� �(��u�N;֋��a-,����O��dU���#��`[Z�YAD{q�bN��B��k����ZC�x�n��x_�]o�q>	���{����Ⱥ�gxc5q��Qjѥ�_2͗��<���?P����[K�,ʴ;|~�0����M���-�z24�>tLfF!G������z^��w��:��X�>�d�Z	f��rN�A���v1�\�C�Z�-H�}��Bm��f+�����k]�h;�-R	�V���K)?)�ͧa�l_���+�`�S19�$�:Oe�Q1���a4�e
Y�p��A�A�QF����p�MD�FP��}R�/��F��a�n����=��p͓���8�F(�ݾ=����G�`$n�i�lu��W��2��kȚWgv��l�:�ɨY�ǐ��YS�Q��O�%-���x��dG�wI��G8#�?�&�#�Z5�-#�N9OA`�k¥��������Sn���,ell�Ewv-�t�oD�A��W袱�θ;���U��
���C��f��o�9��yy�����ߘ�C:�*{��.,[���%��� ��ދ&�-���6N���5ب(>+o����!�� W���Z����C����s��):g���_�f��=��r 	�% g�ٸ��s$)ze�l�G;��s&L��q�*�H	!R�d}�ʫ�7я�ʾJ���N�k3�ҥ��hFTQ����V�z�x����Z����� b~��9�s]��c5���EFū����[���<0��9�g�ܡ�#���1������_������?�+7��n�G�E�#�E���XO7n
_hhK �Z�ݙ^J2������Xb�NC���^i�I���Z���SɁ�09e�v{{�	ˉ��ȫ{�9А.�K�ӌ�V@���-$�M 9Q�����u�h���Qا��+�z#��r\�;���/?�s/�-9�p�ʒ�(��zGi�t�îu.��P]m+�;dCϖ��Xڡ>=����  ����Cx�߾��E������s�~��	�7�>h�l��-���i�[=N�D�eo����y��џ4_fڞ�0U����~coԜ�Rl�S��|�"@Sk1˃JO���#E��dvj���M�D��W��F$n�0�W�z��!VO���Fq`O$� 6�����V���`r�� ���]�qC}�<�,[LR홖~MV����l�
˕�Ě6b�k�H$5� �U!"����G*#�c^������;��d�:�jqmy:;!���!<��S._��?(���m�q�!5�*��yj��7T�]ێ�cA&�@0�KiM��3�Q��[��{��Zw_��Q�6N�dB!���m�I�9�m�n�,&�4�s
����4&�����XS9[��P\�R`�Zq��:����؞�%L��fco_psǙ/֎sO��<�Ϭ�O��D�aEE�:��f��,P����T�c�q�W�뢝�\���u��׼%����8�p��7<Ѥ�����{�洱���Ժ8-�zC�3���ҭ��,���-<��П����;<%�:��T^���s"��m�����Vv�s��2�u%�*��J�|���H�T�������"a^b#9򬴂$v�)}�]f�r�N��@�t}�@��m��g�L��cp����F��Y�{n��#��:��4m���B�����d�G��U�S[!�!�:��<.�1��z#O5 ��e:��õsv1���X��NǓ��'�ۃ�
�tEyy�2x�-��weҾ�Ռ�i񭦄+��s:t��A�ub��J�EK�tO(9�P(0�9&Ce��e����+�؍I���?	��P6�p�P���b�<=���r�1_G��?�����]h!̛%cNT)0�f�soH�8���|���$4H��)�텆���G��m�)��*D�n�i���V c�Qҗ�״�:]~$�_8�}��"�0-@v+x��2,�H0,�M��H4���&�����w֟!:S�:���B�Vw[����Glv����3�_���/�A��G���狹l��Εթf����RW*�qV;�{������}���Y��ܷ�Y����ᴨ-1?�=�Or�b�l�?K�����A,r��u{�<��=�B����:)2�^֠r��9�ѱ"{(�ރ�>PQ����/O��@����v|a¶+��Z����~f��K�\��4=�h�ӝ�;ߋ����f�YeH��ץT/����z��m�m���]LLF�b���I��#/���^
IG��Ge��Z�e��J��6�'�U��<Eٝ���~E��+���k�R������pMHfF� ��K'�N��o�G<gπZ`*�����"t�CH3
kUQ)P�~��L*�Y�e��V��|$P��R�� �}~n�	�^�;z��)$O���Jr`��Y9eM>Fx{(o��1������Lq��Ќy��f�Up��$��fz��{Kn-H|�ޓ��6p�'�����f���KP�+㴰�w�tZ*��3SE�'�?Ӥqk[>q�u#.]9ǢFD��U���N�����/w(�B
�џ�`.�@b)�M�����(%i;�^�γq�X��IJ�O�%1z�x��p�^���1J�S�8������u��k��Gcb��T�Ԋ�M�Wx!�W�e����B�u\	X
�w��U�_xwnB}�@YQ+�<��x�%NdR��Ǚ��f�@dO���Ds�Բ�.5��i��/F1f)��P~�j.�1����uW� ��Df��hxq�C�MH��!.?�����T��h�6 Q��$N0-��~=;�(�� |�ۑ��$�41�c+QŴ�$��)�|�h�#,q�!�����!	��D��`�eQ�� @�Є����en&����Ƅ��Cf�gթ�#[�b?B}�J ����,W��E�$q�S�k�rpl�_&@���`��Z04���V���GY������&/ĕT�c��	�����u�K��YZ*��`���Y���<�Cg��^�ަ�yEX��j�,A@�V~1�����D9C��ʀ�"���"F��H#������j�-"�u�X��Ȧm��Ԧ\�'CDG��N�]�N����i�X����W\P�PZ�� �fue�F��w \��a�\ֳt����)�� H�\�#6��o�ǟ?����d����;Mç��s{�����e�C{�Q���s���gJU�&lh�~3��O�ɱ'����}Ÿ�D�o��u�Zo{��a}(�G����Bo���0R]UQi#��F�ڀ!�E�e�y8�e�3N����.�5k�B��vy�6h�KN�OH`G犐/4�u{\�����}u���z�C�����4HD��įq�I�*��\̜4�I� ���34nu�?c(w��	}�7»O�'K�`�p��$u��YP���K�������D4��k~]4_�UE:6R�6�j�0�D�W�Z�;a��o����6
�������%��C��S\C���g�3�.pJT":��	yo�sp�&(�h��@�����Xƴ@V,�����{��bFQ��Kݐ���}�GU��Mb����T��za`��fOZ:9*�A��5�V����H��%��LuY����d�6Xî��k/�B;Qxi8mȑ0M:^o�$�Dq�DC8P�M!�����H��#?�"#��w���O�֭�j��ot�����z ^<	_�]~m(N/�{���Y�^��rS�
G=N!4���o%���M���[�=�~���	b<��/���6n���s�H���3B���QX��)��g� 2�[O�LVI�}�T�7y4�TWL�bIg�o��3�OP�o��-o侇����$&ü��g����hx}A�8nYk"��v�a�#�Oi�Ӈ&�9
NS�]'��g����1���Y6qz��Y���j����~23 ���pn�zE ��^5Y&�������1��/�E�'?��TsuD��,y"ܣ#�Sz�o�Po��_�U�2�~%�=&2�-�?U��ұˍNjZ��R�j�E<S	��V����S�W�?���E�h�se��L��c�xL_��EO��Fj�)���(�E8d��I>L{�2�������-�v���	��?]rJ���~o��xU������Ҭ멒@WQȗ�%��)��V�f�*8om��]Z}��~��[VCt�n�
}�Ͱ��Z��\��a(K`Ւ_d��d�i�ޘ���\� �<��C�j�\��l��Y�"��=N^�ܤ�0��0�
�՘�ܓ%��W4]~Wv��ތ@�Z��?���+r�5��iUJU��Y�p
S�05ȘܫIhS�Y�"��hu^I�-)���f3BR�n��d Ա'�������Cj[�|G])�e��V?-hk q8Wŝӟ8�D������nUx}�l�.�R��O˻:�.1M�"��B��� fa�&��-x��>>S1?��q�w�C"���!���h(90��a4K�5��I��')�c�r�tr+����ւ�%D��Wڹ�|p�s�d����A���Ϣp����V�E��V���\�V��x�0�]���w�����oi�CΑ���BwUD� �1���jRF¶�>'�L��R��v��5����J=z0�?�����4c��+�:GDuE4��M/=����&q����T�j�>��ؒ��·�/f(E��9�"A=�b����.qn[�ำ�:W��"�B𑠓=V=�����cr�[;���G��?�&V:��M
���)F@�|�/��q�r�����p/� e,��mI�h#5{�H�ʺ�9n>���<-�9�����W���D��(��4;�V>� ��d�ȱs/�H�X�}����
���#�+7�2Ǫ���z�h�V�K����>�o����&��}�.�%>�n{^\`�|�� ��W��ۈ�, Ǔ!�si���f
<����7���qn`��U��j�,�U�ӆ�=V�'�Č�z�<M^O#5�F%�}ʏ^_9��DT�|L-�[�!ua	��� ���K2��+lA��� t���(>��`�v%1zZ*�m����V8�6ȱ�,���<�->�k�pf��Pщ�Ȃ�
2����p��zV���%iM�R������Fp]�Ư���0�ѨE�V�r�����*��"��k��$ &s�!�����LJ4сi��|��E���%\M˅��� �@T�zU^P��;���A����q&�:�5���oRkOs+�x}\n}l&  ��N1޸�t3N)e��r�'fh^ʹ.?�~r�	�1���^c��z�3��[�M�0)���l���hx|,�(? �C���נ2@Xca>�Yj�,y�l�X/O��1ӂ�j����%�0~}vZ��(/�	��7�z-�g���(��]�=(��,Y�-�y\���&�)��X͠��яť��r����!+��
��v�B����u��S�m��Ji���t�n�Zi�y��j)rƈ�?��-[�?kF��1��G��ʎ9�Xk&���2��Lv�A��xR���F�Szn(Y�ŀ�2�X%����t8���\�rywCq2cFp�<jϟh��@`-���v��@dςBm	�\~F1�^��c�_\9�̿�BuRI���s}��9��6�m�'K��PG�wF;^=4�m�A^Z�Eu�
MKe��O��vcB�@�ER������6��;���7�ʂ�N�s�h ��w�#�B
�~#��������
%��
�P�}��ޏ�����Gb(�$ D�|K�@l^+����:�-�B�N�!b���Ot����~�~�U�"�f��nS�[��qP*L�y���߆����U�s{K}�.^B�S ��<�etgE�T`v���Ա�kH��eDŃiw��v��*����Ojc�y��/�7X��,���(��hw�'f5�ɒ�ǜ��aGHT�N��#�:��]��D�it�+K�6ӆ�6�HQ�}�A�7Õ��F1sݦ,_�d����]T�������"W��G�����-�����F�}GC���t�����U�," ��8��ZO��
\O\Rl��}��Ekwn��Ni�;��;oAI�ٗC�Ɂ`���N*�!�A'ؑ�u��C�brM��/��O��t9I܄�!�Hs�jN�f���v|��Y���J��UZ�C�����4���������ِ��l��
�W`0|Tণ�`�3Y�ȿc�m��>���	�͢�(2��dl�Cȓ0@�)T���2){.Ϥ�߻E��; �[�s�����6:�T+��R#�YeZ�r�*��=m`���A����ۇ�6�m�_r-�a�,�a���L5��Q��J����֥%�}ޢV�76��7߲�<F_ڐ[����wo����[����R�("�H2��l�H���k��r��(mV��������W��������rjf�bR��RO�X���Ђ�;�JVu=��z����U���iJ� 6�{�O�X�l���j����=��q;0q/��Ѯ*Ζ�۞��_�̈́G����5o|z�n� MT��F9ү��m��c/SL��RXTV2�Ó��m������ q�[��bO�t�����Q�_x���+����S���e4̹ja�"�l��@7�ȗ����s�$ڼ\�K�e��6��)X�	�S߆i�|����.���	�eL;"��6��'Iy;�GLR}�Z�w���9��b���[W�̡3�e_�^���ѿ�]�{�uwĴgx,�S	�˦���^�E@�IE���8ؽV���Ij��������,���Zc#�~�Ke;���}�Jn&�=_���-#T�>�Y��ȳ@� ʿ^�r���ş��}t��|H訵�svf%���F����$w�]�&~����a%�"�" �4���Zf�2����e~�p�q�麊��+4���:,�#[g[�~�e�ˋ:n͌2f��1Ґ�������C���%��~��B�8���,"�$�xy�o�~e���4`�oǇp���a�u_�u�2����"�h�ˍ�.