��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��,�y�}�ǰ�=4d�H���`I"��W�`r���T:tB�T4D�m�)�	1��I�t��
��8(�8t>s)ו�."[�漆���]�~�]��;�O(1#5�-� 偙O��QZ��~rL'�x[�i,mׇp���O�I43��4d�,�H�����SN��d���3���r��m���̨T�I;uj2Y� Er�*p�Q$Gm���p�V�`�2^���,hz�<p��l�Bxt�5��s��\yq���#�@W���f:m��T�	,*�񞭋����_��㧋l�	�\�:��uGd��PǷ��N�I��_����Tuv� ���us�(H�~�{2H�:Zor�Q	#%�3ˠ!��iS��95�,?�.���/�F�i{#���Tp5����Ҥ0{%���2vpn���X�����@l����3dc�ק�3	�Ed&3�ZN O���z��s�yxӡt��v*}ԫy nj#��lc��m戭k[��5)�A#�����8�!�]�Z�s�M���t��w�!��'ÒE�rv��Ϝ�c@<U��\tq+��&|�&X1)C�����r�A~��B�&�����s�:n{p��͠R�X⺂L^��R����c���f��J^?��ܣR�O 1�rV���:��T�4���AD����˩�F�w��)Dm�O�b,�a���1$��c��7t[i2>�ޔ0,S���󧇳Ϟ�ᒨ�-��}�!6��Jyv�醊�^_�(�H�(y^����o#����X��3-�k\8�M�T�"`R�DF6ȕ� �,5�;Ҭ C�k���1\������k�t־9�}���� ���QHF��"��t�9 ?��{E_�7��!����]���-�p^8�3 ��TLM��q�"��z�����`%F�zU��K�^�Y;FI�$�*,���!���w~D�A�]�#����u/��eס�yl:TJ�a�ȆJ?fgu��!0m�e�ӵ�:*���"GH!՝^�"VIk,P�;�Lۃ���Cّ���F�O!�
+y�Os̕��K��u#���dNh�/��HZ�=�(G�f�Ņ$�/�Uw6��@nK��q���*  ����>(��x\})*��耳K)��e4��3n��zR��^�y�&�Q�`<��o��R��.�$��`�b���UM�ˌN�}ťH{�s��&��y��.aW�E���2� ���v�ˌrr-���/�v��
��R�.Z��@s�� ���_��'<ź�}N���i�1���P( ����G�&嶩�{�d[=�~�F6	��oP�]��g�U��Ѹ<a�|X�Z���7�l�-�n*�41>�2���#�ÖZ���6�!3S��&��"r�I���0W0i<����r6���g��"�Gq�`XK8M��y�
��b��@CJ4�07�;�a밽%���|�S17h�9���8C���܎aN�5ឣ��������r`0Ž�������"���h��D����K��j��ԙ�y����K��ʫzA~PYFȦ����#g't=[�׿���S�4a��r�@���Z�{���w%TE�ef[�$���� ;~��G�¸&H�OD�U� � ���\&�L4�/�^	����w��u�=�'��w9�%�c_�k�X{[ ^��m�����ЧI������,hJ�'�1�E��Z�&)�A-��)��Iq��<�ω��Rn+�:6Z��Y@�8^m}M��eS���lg���~��'5�|�9�n��3��&��Z,z�2 8����ʳ���������{˵y4�_���j�=��Xz.���LNV�ף"CNn%�z�߅C�� 0�4�z���X^�sV��0 i����uʈ��*]��7��os��{#X�
	H�$��]���M�95�6%X���3}��|f�$A�H�J[W� ��Ϧ�"w-�1�������Ǿ�۽�^Ws��8yͫF{�PY~�¥'WXp���T��0.0�h��	NRS�BS�7�ᏻ����UH����j���D���?ׂ�M�)��2�0�m��X`\�ta.��<���C��7�@yW����$C�~@zq�=#��??��zF#*�`+^�u@P2�<���u���y����v�<�!�����K��TH9H��*w�G��M���"�b�Z}�]ݟ�6��pN�t�!BR� ������%O�����i�i����R��#�~�n�뀽�%_{���\vh�#�����1�_0"�����j��=	��#�ĭ����"t�����(=4/�Xr��[�5s�vF��=)/�/e3��1@Xqm������J��;�d�e�_�6ۿ����f\�D912[2)ނ��L��o�.涑�������G���D@�*�t�t��R(�XR�vN�v�U�뭪(TM�ɖ6Na��B�\�R�!AMT��E�h�q���t�6�^��2�$�rL�.�����ۗ:>S�є��
�]�T�]�uȻG	@����/�O��k�w�!��+��Cӥ�|I$���@'p�c�֐�g�r@��I;K^��zr�ˊ�