-- (C) 2001-2016 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
BwDFSaM1MCAETBrntPX0Ob/q2JhlToAoZPLA96EPmuDi07mLl1CJYYHi+N3Cc+K2pqgNOtstwqQ/
oixoM+eDRhxwPJ8mUzrLyEEAazky2vb4SpuFivWqITyRFr3AZFOKtqdCmdLNIIp67pZ/560I1sSG
IdtKxZ53vAtDPPsEQ9xi4EOjMSnSokNCO8f4rWUePkUFFfVKfz9EmApMgMIDJ/lfqNyiiFp+cMOp
kiojHpsFSiHK4eZjfzMvdT5tEpJtxwI9HOGjv+pYFKXMQkxxy+U0PYREu4xC8vGF40rQIDth8ToE
mrkaTolN1ncteVpaq3W1dKbLBoWN6SqEjFd5yA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 2576)
`protect data_block
ALZsDik2aHCp4u9OUG1qH7RbUQmwl2EQsWIZLlIhEcNc7ds2zmBXyQ7lUpldtLvH0Y+w/kTaAtBo
pHapuYShPny55hhiBhsNBvwE3iH4hJH4sMG/N84Oc3XP6xRgADndkCCjzTvbszu9pJqqfKFPEI2c
mPO3pBAD6tTJ+s5Z1++h85WYDAIO5a4mzoddJwscXVAMee/T/eyjzk8tgTF5vXMbdHRMPob9y2mT
s6jJ3FYFHvr+fTmET6X4e+ZHicvNDiarATg224Ofxe1kGAGXFD+DYXIOmHzr2iqBqAQdmLt15DCE
Sku4vK5DoO5H+vuuPSfWz/R2e+9gaiOzOPHaUsxql7LDzaJhLMEGO8yET9wlbTAYUKOFspa+Z7oa
B37Eqn7+BJ9p3HgyMESTW04r2F1LJ4371gixP35DwCnR9t8CUoPOGOQzkPSN534+/iagTowp1i30
n4Reomnl8IW56BxufGb/F7e2iSVn/3RaJgXGMBuwksYiBs3fmFEX3qGG3aD6RYAyaDq7JBnUHmkQ
/HNjbIfHd2nLj00zLaCIcg23blTy/UtisWzaf8Rqlq5fDX5bqumZmqZhnCyowpkbd+bionjmFPdY
oYfv5Hp8KPOwuDSvybMYlTTx+D0nIOBxpd2dPBkFOxz2BB/ITA48tlEg+8NjGHNRasr6NBFTFaqn
i0TyU6vBaTNSCcAdirriXcXDpfWaQPbbD8YciRIzKuWXIiNMRMSavDQtOlCyiN00u1EbgBaBRZ9S
uwngA2VanxYSsYRWZ9CgchGgGj7OP2CrkuSrOPLuKf1leowSM42VAvUU6BRwcNNbSB9clRdS/K8j
geKo6CCL56mVXF1EU0U70luFo7lbiP3zn30BBkIwJePi+IfCg9ZCDPR8Ky8iWpwBuD/OxReilAIo
vTDg1tway2YH8MKRGiUqkso7Kaq5vJNn+G0CFwJbcgw0Cs8Re6A6Xqri/+2Hi6Q/nM6pT+JqgGy+
Qa58h42BdACjDE0efuTyS2j+wIuHKNOJR5OXsvks5FwdqMKV3+8vPF3a4GlgU+FU042YVMyb82Vj
OcbUnpcOnM8pk3AszBZ35JqOc1qgN0unU3XBH/dHSK8FUu6/zBUX3OQEdkthoqGUGfjk29C4h3gi
crMhqne3+wqonk24m52hoSfgV4lmCRAgLjVFb5xqvGsyC1BOi45JJiz9rBER2GF7ZJkSrojjm0ku
tVahzc1lKi2cVkUUMItsXTdHe1WA0p9uapeomdfs4fwvkQrkTYWBcM+z5TAKMxk1xtVmd+Erjcn3
H528LXketE8ZB4kZ1L0pHV80SZ42NLhHrkjDnQ03Hdf+280o9xZJcMUP8lQzaIERMJgHAa87RrBo
5rBmZdw4Otk2K91wcQyq1iTS/D+A7zeMWYKRCxfY2V/BQp3ZkjMaeU/8jAKep3I1J3NkrkEaJy7Z
qpRr798As5F81mM36EEXtzYSvGmgHgBTU/yLSWKnPada6jAHvo7LgIoNVW7TbDL+P4jnzbn3c2uj
iOB5u2jYxUvrVbhiP+vp4EuicpqsDARSPKTFWbKdsyKfKttk7PAubh9Y/qxXoEvh2+ktqRBtScqb
NRrTu0KRMmgdrC7GP8LyXRxmMZVPrw49X6B5a8PBwfgwEeTeLMKI4xdROYnBMVQWTF+HJWLtdC41
4ZqI8MmFEJxu7iLt3vXj1DzlaOJ5J/D3Ry+caGybqxp/h3og2c6pOADF1Lhg6chfQ8v/doodPFkl
GUYBfyTlhvRr+Qzo/sMsIHWeBvRT8i0EM4oSJttMyLEI0CtwwMObn7eD8V2c/80/k8BvoRERVGyO
FbV5bwe1z+fRXXlo1tsKIPWsMcNeAIygyUDD2EbV0pU2jd0P7iZIS/NoZlt+MAWy3dAFByID9csf
lAvyBrFRRLj7HUzn1MSlnrnPw+l1pDOyqSy2Iws7sF5yNJHOql8YaO5AzhWPIsINXC5x2aYwLtYm
0/y4UDVmOiSaJlOLBwLjf3QfUX0vUWPqiLRVThyTJqSFGQE2dKainvjvlAnTBYk1zOcIV/ly8lxS
98HWzE0GwHjURmVaHNR9XatVTJGoGejzWDGKu46sKK5wmmg7WB4nxQYvMFCAt7KP+s2jpVVnrbTy
b+kUXUFiqhb0aGuNSvNTfgm4XQzoxmBqTrxAHpNd6xiFATt+yp2JCkuuGEfX75gGMcFxzI7GHIpM
t5uF1dvzqLC4AxTpYN01K6HA1yBP61+ZWgELuhUFf4BkIl1NScQn1ax8JciZt1O++enIv26TvMNx
XqDoOny37Yrb8Pzem2dnyJBJrZNxr8L01vWR8QtQ9zZyCPWsfWL4gIAsJzO9VjYWOauugo9W+zYn
xlfKGWeFkmb3AyES33lIhnsURy5ajoxxWwF7BeGqkpaim63rtSNyktc/I3ykfXggbs02axu7siA6
8KYTDPbj/pX84Ia6WWd/qEVaVYjWfQ4k48fSqZJPkzi7RcONnw9BY1/AVIUwUOXpB9m40us5Y1iv
aG2uGzetug2/AHZ/dfhfbr5KTkqIoWgdIdAK5nOtbVO6tLEPgT9LCcRv7a5hoTbQjcG/MSvhaLcV
awz8eb9VCe+yPM1//L7VN4MxXjFDDmB9Cq38CDo9o96riJaxn9LVC6nJ/Q7xJEK74D0I09X+GA6h
LbAWiky3l5t+3HxPXDaYNEO7wIC0jp8Jxe/RXOb3eIowk9ZmqKKVWRoAvvuuQajx1mDty++O36vj
2beE4PMeFAG5NFseKQ/jgBT+zrb577083zmKCV4IxrLThHSLc1FecBeO0SoO0YrY20IM+sFka8ks
4xyZFiKScwK4TrsFloP3eAdFXXELFTvHr4WlZtBlTleCNYlu1Kle74M8C+t9mZq5cddn0XNcjB0U
AMPnlk5PEHCI/SF66GKY+veIR+d9NJKSGcFXpGQ7iak0MF4d9mTTaJpHBUa1urpf5IdZJZoYbWnv
b3tKvgcL8YUeaPix3XaGQPE7EB+EJDAYXQDEPITPrMZlVnhTTzwau1zYhy+9b0ZEPGZ9pcj2FXRZ
FpNgcwDrtVzfMBp0Jun0AnS9BrtFRx2nRa3iX2K8aGYLFqHiBZ9e+C/xdYTdCOx3MisRBep4He3x
/A0fh3ZFGcnCMpKi3MxCVRaDg9RkBNDi9SNksKHibNpES8lgBT1PigbWkKAjGwDqReY+YZ3Tl4at
SJ9hCqOmmJlu4Ie5YBVaZ2nZsUVKw3aikJEhxEuPk5UFpBpg0ACw2XccAJlOkIbq8QVsoEYYtK3z
6tKBeFyKUuygvTV5YzoDzzkUknCz395ro8JILUw58/+0W7ZQiAj+1fykzkxhg9/LRnscEDJAeRF6
c58z3mnYoFpxVAW6NdXsnPzL0/ff+tlB49eOdGEbTxO4PY6yC21C6rhcbem7METXemGi6+wgyg2/
q96KKE89bK0sdt8=
`protect end_protected
