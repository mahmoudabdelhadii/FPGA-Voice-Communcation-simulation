��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����N~@#�k�0!����+��=L���0�ԴZ�2�Mc���ZO�����=�����վ�	"cqw��a��TS[��{=:�����K��-�մ�(��k��N�-� 偙O��QZ��~rL'�x[�i,mׇp���O�I43��4d�,�H�����SN��d���3���r��m���̨T�I;uj2Y� Er�*p�Q$Gm���p�V�`�2^���,hz�<p��l�Bxt�5��s��\yq���#�@W���f:m��T�	,*�񞭋����_��㧋l�	�\�:��uGd��PǷ��N�I��_����Tuv� ���us�(H�~�{2H�:Zor�Q	#%�3ˠ!��iS��95�,?�.���/�F�i{#���Tp5����Ҥ0{%���2vpn���X�����@l����3dc�ק�3	�Ed&3�ZN O���z��s�yxӡt��v*}ԫy nj#��lc��m戭k[��5)�A#�����8�!�]�Z�s�M���t��w�!��'ÒE�rv��Ϝ�c@<U��\tq+��&|�&X1)C�����r�A~��B�&�����s�:n{p��͠R�X⺂L^��R����c���f��J^?��ܣR�O 1�rV���:��T�4���AD����˩�F�w��)Dm�O�b,�a���1$��c��7t[i2>�ޔ0,S���󧇳Ϟ�ᒨ�-��}�!6��Jyv�醊�^_�(�H�(y^����o#����X��3-�k\8�M�T�"`R�DF6ȕ� �,5�;Ҭ C�k���1\������k�t־9�}���� ���QHF��"��t�9 ?��{E_�7��!����](�S��0�q��w�9��=�i]�1�GʦȪc�W�XC�|�$��}q�6����zf(����լml�dz������*�eLD�*�,�m�]ہ6����D�Gw� �g��' A���FX��\өܹ&�6�h�Ð�$�(+��埧��= Eza ��찠pr[�c&��nP��x�2�TK�M�V���3Y4vIR\������ɭ�1՟?4�_y�y+����ƄJMm�����*�\F�Z�� �4�Ϩ��8��$�A�t�- ;z:�̌sA�w�Ħ�J+�꺲/��r�a�ΤO���x-��~L��QpXwKC�T���b2^����&�IJt�`�������J���*2�vr'�w+e�ǩ�܈�0�2K���@��8�|w�����y��`�B�4�r�7%�]v�������ѧr'��gHD�)���|^�ėm�/\
�p����"��9��(#����&η�ҌC�J�e䒌.���y����L��iRx�A������"9U�'��b B�mZ��0�~Z������q�f7�w2M;�h�_X�7_B��@ �>�X��@�)e��>�#�N�^���o���'��"]�݇��Q�܉�N1����<�`�B�0C,Q<T�+�ƿ'eM���/-k�.���MJGx�{z�͖>"��?D��Y�� �l�̟r���)}7�������˗f�핂HE/j�~ȃ�b���ՙhU�y��x��G]k�<�hƎMTcLk�.�Qcgu�6��ʾwe �gk�&��B�h����]!�N0;��R*�>���\���MSt��1���X��˩�8�?�YeY�$朗ɕ�Pn������Y�6��K�`0Ђ�|��Ҝ�U�`� �K�V�@�}�`�N���/5���1�{X�}x���Ȕj��|�M�.c@�:xG��Ȧ	�VW
�+$lmvh��#Gd�F�a]��mp��1�y$���lB��J��++��q���E!Ə ����B����q���9��~�^�J{�=���_��5?E���YOv��s0}�m�)���r	0� $�1�mM��I����2:���&A� +�!R!��O��!�j�F�A~���1�������3�)�'E3��O@�����J�R`VC	R�0ɮ�D�~�f<�w�i�@�tأ�:�/q�*;M����!����g�����!3"d��M=���T���}PF9Q$���O��⤍2;�8g�Җ�"�+�%�IK�[?51���F! |��NOS����4�1��.� E��`d��w XD���܇8�2FpO���j`V)���F�gF����΋x�g��`q���E)U�KǨXކ�Lp�$ϵ�}�r�i�W��W\�-p�U)Q�0ftp-1��.ND�mv��rp\a�e�D�ٟ�b?��49D�O>ȟ$�F�N�'ᎄr���g��/��Y��{�EQ	�*>�G.|(mtVڏ=���ȋ�$���%ZW���Q�jP�۲�?�	~É8ك�+��yWA��q�=C�����+��J��5Mr;���e���帉�'�V>��W��6�`�;R�K���\����ʊ�o�� �ݫR�^Բ��
̟��]Ks/X\���d2*/��/���QT��B;�-�&Kv��yn��.���6{j�������/�2�y��j-	{U��d~����l�ِ,Nj��c�E��"e�q�
2��m?L�k�����/v�s�κ=J�����Xv�Ox#qՏɃ7�`��A��f�&^��+"�@L�W����8�&�� z�G̸H�D=�������`�~�V)֡nα�/k�K�<MS7��W�_�����N]f
��$������fy�X�Q����8��P=��O�͆�Pn�kƣG.�;���y�L��X��a6�m5�Х���r�{�h[�1L��8�	�`��g�hz�sU��?�k|a�fb`�8t�\[,�
U��5-3�ʗ\�׭�J�h�3F