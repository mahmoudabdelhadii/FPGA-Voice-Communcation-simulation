��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��,�y�}�ǰ�=4d�H���`I"��W�`r���T:tB�T4D�m�)�	1��I�t��
��8(�8t>s)ו�."[�漆���]�~�]��;�O(1#5�-� 偙O��QZ��~rL'�x[�i,mׇp���O�I43��4d�,�H�����SN��d���3���r��m���̨T�I;uj2Y� Er�*p�Q$Gm���p�V�`�2^���,hz�<p��l�Bxt�5��s��\yq���#�@W���f:m��T�	,*�񞭋����_��㧋l�	�\�:��uGd��PǷ��N�I��_����Tuv� ���us�(H�~�{2H�:Zor�Q	#%�3ˠ!��iS��95�,?�.���/�F�i{#���Tp5����Ҥ0{%���2vpn���X�����@l����3dc�ק�3	�Ed&3�ZN O���z��s�yxӡt��v*}ԫy nj#��lc��m戭k[��5)�A#�����8�!�]�Z�s�M���t��w�!��'ÒE�rv��Ϝ�c@<U��\tq+��&|�&X1)C�����r�A~��B�&�����s�:n{p��͠R�X⺂L^��R����c���f��J^?��ܣR�O 1�rV���:��T�4���AD����˩�F�w��)Dm�O�b,�a���1$��c��7t[i2>�ޔ0,S���󧇳Ϟ�ᒨ�-��}�!6��Jyv�醊�^_�(�H�(y^����o#����X��3-�k\8�M�T�"`R�DF6ȕ� �,5�;Ҭ C�k���1\������k�t־9�}���� ���QHF��"��t�9 ?��{E_�7��!����](�S��0�q��w�9��=�i]�1�GʦȪc�W�XC�|�$��}q�6����zf(����լml�dz������*�eLD�*�,�m�]ہ6����D�Gw� �g��' A��)�m���b��ӎ���o�6ūvO��=�W�������}��	����z
��z�&�P�K#�^Qץ�_������&�)�ٺ�u#uD�	' �/|�qf�M&P)�tL�x�?�u�����ҽ�����*c"q/�\��YDl2n֢�vtX��Q������ǰ�6K�gVL��ο��Q�������-�˚e��"gb�_� L01�D��ثU�8-��Nw�@�$[�>V,���6�����=����{>G6��v�����φ+Y��	�d�A��b<�)��Gp���k�(�vWu����!5��YB� 4��
��<3ܹw���xǄ�'����160���C�sA��d��K>C��<Q����y����d�p�V��5V��ά�hTR�qX��vW~0o�[y)�H�����1�a,B��f�(���b\�M5�����E#އK��wf�b��2�c�OA$��Qhb�.F<��/p���o#�)�٥��R�_�#tI`����Q��gj��S-9|̔WT��b�$�f
��<���*$a&�'~�]A[�>���;qW�Ϯ���N�+�\2�x�tS��OhT�}�m�+O*�&�i(9qجV;�kw���<�D,����`=�'�[X��<J����(;cL����R��3"�[�j�zY~�sX��w���|��^ĉ�V�����˔0�ٍ	`kDڲO�>���4��3�^����R"&��˱�'�Z���a7�D��c`QLn��#!�nY��i0��y:�����)Z�S��� ��$�D�w}�1�<�����]^�q<�����qQ��u��z��o�T�V���G�6|C�;��0c�*�o`��M�2�a"ǐ@w/ʝ�����sK��A����*�}M��4�$���J#�f���`1Nl���م�;��B �|��[�)�����ַ祙"'���Z�͸�歵�>.	-�B5:�����ɕ/r��]M�U\�.�|�|����$�jv�d���i�6��U�5��C����/g�!�OV��9�r���*|3��iڂ{���T
@�
CX�Ͼ�@!�{Fg>�����լڢHg	!W�S"*"}�*��}�n��r,wb/�.��tI9h���e���-l�����8Y��	���Z�?lN������:���&D�qb���9��p��i�9� ҝG}Ǆ�{�-�	o���k��79R���9�0��?���Xî7f��Cfڟp�Щ�&{P�[@���؍���AqIj��&���[�C0ݍ4c:�vd@�I]"G�Ԟ	��jme�Ga�>bXa		��{��&���$(�����ͺ ��f�HDƿ=���P�� uA<��Г��}���=���ƥ��za�6��n(���(��I]����vB!e������S �ESbF�g�C�[P��0Z��(GPq��U*���-,�To]"M�uG��S���#�[y�J����S���B�ۖQnť�iWfcK��94�D�F+ӈhf�G��
x���g17�@t�Jd!�	:��=��Pd�F'u�ʎr$��Q��v�N��"��u�E�N���$ѯ�b%��H��5�CDwR�tc����߸�c�;7�a�Vy�/��fO)�t������S"�&�}��?"�ͺ�08�~�?��=.���w~�::c�B�fvnv���]4b'�?�f�-Ke����%܎D�^��,���
7�Ņ����^+���mK��#��M��9a���0c^B0�vO�Y#��h(�"�:m�q|z�h�t�]��Q�X��U���^$�/��W1�#:x?�wq�ŵ�!�}��G�ZOu	�
Ҫ@�E9���A��u��?����C�\�]�}��6�x�
��I4�<�3����e�g��2�]�)))RhD�
���Kw�I�b��e�@�e�n5������E�hG�H`�]�k����~8}^ChRӺ�G)5|���y�׍jc��l~�مy�)`�!ہ��'���|Sܘ󬰬.���1��s��%��#xD	A�ܩ+�qƯ�U4
��� �ۺN��@V_�c��%@Q������F����;���]
�d��8@������
M[=�e�R|a����o� �:nT> �YX���Uq����N�jݑ�|۞��s���X�\L�h��b�w���ԙa�zu��//�x5�мz��/���qb7��?��6�3.<\-��CX�����:��P���{5�B� ��䕊��3��v�XG.���E�	>P�͇�'��w���0m� j����)�6� z7*T�O�AEo�0{ܨ�z���AO��P���� JK������ӿ�6��# '˦�ys56;k�%%�}/�����/}i�{�=ʛ��_�x� M�t"l�P	����'��9pd�|[%~ʟ�o����7
aA�]پ��ړ�u�K�M��0�ɞ�����;B�Qc�Ֆ��{X�s=Y�����u	�m[�uJ]  $h�F�aX��OKN!����ǵ��3 ��$V"�ĭ1o�.��\�7��}!Q�	�����X��]���L��S�������|��$RuH���!�9BE8<^o;Ȋ)��C+��vs�Z��]V���f��5���M�
4dO`S
�7,)�����3��m}$0�����z�u5˖7N��`��/��,B}%�\���&�I��E3��A�i%9�7�4p7��փ��@���7��f��K���p��!2N�s@�hL�= �+����Lt��/�v�� $�S��\�����6�a��!v@�K���;ȡ���\�� ��=��L�H�����J�;�y_���St zLF6��h�n{�8�1��Rm�8R�3>���ivt����9*�d�|�{���HN�K�>|��B�k�_6�䞻���<�t�
 ���+�T=3I�4��Psa�RWi>�+45�/Fɚ��e#M�	��_io=�<�a�-�����AG��JF=�i�J�4'<OE�!e9_3X%1�6�ئ�k@={_W.cd�{�?V�p:�PU�	�x3�۶K%�nc$�u������I��ڗ���ط؉���_�7�Sx�ұ�c���'��y����}��^�ſ��)`#�ģ�G�^�����k�y"�F�#QsX��t[>�pQ=�].�B��S������Y�����d-I�^j�Gq8?�l\GM f��Z��@1��Y����v�}47�P{��Ȗ��S�~���]�[��o���a2Z5;W���F�3N�Rm�ڻ�{d��VZ��x�`j������$�ef�f;�[��U�S�V];���b!N�څ�)���[#�9��>~�Om(6�Q�)��ٶ ^w�7t��!�@-Q��GB"~�Y�����"���F��qu~�"r+�47Ս�+�km��̀d�/�:�|��d�<�G�d�Ⱦvv@MPɬ��,��{�r��&�r601��j���dp�OŲr����!Z<L�d6�R������8�»�V$NG\?�ͲS{ܛ	���4js�/6��V��;0]R�(L���Hd5�T��{c�A�O5��JS�k�u�ց�r�iI�y���K,�A���F���,@�Q//:]:m �SarI�^��>�2���bx����@d�b�m���<SIx~�#���j�����eh������`>T.)"�,��/��F�S��=��$A�����jk;x���Gd���7w�#]�M7s���%�řpN�	����O�K4��T��w����$T��5(�Y��^���8ގ_ǖ��Z������V�6����o?W�h���h&��CH�g��i��cN��xRTʒF+m���9'&�"6���V��w|Y}'�6�R�Bx���A�1�Մ�+[Ng��=�8Te��J�P{Y�مh�u��֒!��������e�$�4�b���곂J�UN>r{h�SV'^�����3O����3��h$6j��xT��i���ĔïSi�r&D�pGm/@IF���{Z&�F�yE����Ҿ�k�I`J��	F�g1v���ti��7����O���#Ske�d���x�lBOOM��������L
Aѳ֧�0��1��7�	�B�`n����ᨪ�YpZ�d��sh�b�w���'�*���8v��e���m�ɪ����8's1�&3��q��p'�'�x�����-�Ѹ9*�	I�b�伫����]��W}Z?՜M���5@���Y�A�od҆��W�M�{�2��R�4�аa�ݚ ć�d�`9D���5Z�CK�~n��Wq#��\�ƆM/��`t�?!���~m���x.E`l���cE1�:���	�8eZK�݋���7m/Ū�T��Ǉ��1����&�׉�(e��‼"��Qk���O���5
�P�0�uff���A����~_��u���m�l"2�L9/������u'��	��a��⯋�i*��r�Csj�� v�QA�C���e%'��� ����P������iEIY�tA��25�Tc:��7�'���*�����٧Ѫ^�)����һ�3!G@D�0�睒IM���;I��ܡ�cܔ�Mش�(+*�j�񝯁�@ܓl����P�N�Qz;6�����hLhj��OW�F���}|j�M\a��<�|9~ч���rb$�����h=Gqˀ1�����ጣ�N��p�
u���j�$��h����Jk�k�טSֱ��K�o���M�8�@Eﶇށ~����-m���Ctx����z�%��P+�`�]dD7����?��MF4Z9�]b]��(��P��Q�jc� 7����i�b=Y���}�-�}��/+O�!&a|\y���8Wz|������䏅mF��~��8�A�/���ڏ�k��R�"�TW	ܝѻNŨ!�(&O>�2�=�?�p�X���W&n����5*Ƿ��{�p�\u:Df�s�Z�-�^`h�M���#�)���;+H�.1qz� O'$�}
��l5��g�,鋄���Jk�1L�-�vf�(P�C��4yi;-i�CJ��k�������`o��A*H���jZ�����<Zm"���*��Թ�����vӻ�cC���L	�k@�m\�K��|}_�f�ߑ�0<a�
u�?3�_����A�F��W��fcӭ��x�7��S�xfUJ�ʙ��M�o�I��β�6�hw<~���d�fht-hG�1�6X-��Ȳ�Q�-y!�R�m>�J��#$T�T�q��~��&�q��QBC�{�Tc(-�f�`n��u��qw�7��tm�8�Å�xP%��v�s�F�>0m k՗��j�eEEv�͍����943G���L�H������_���_ͭ���Î�xC�e$;�D��FoK-�ЗL���
�WC9�AoZQ�i�?�Y+9GE�	m� A�iӒfv�a �(a/�-�K/�`��w���)����ѝ<�؁�~��o�L�a�1�FwVȄy�Y�4�^jw$`S�~�m�}��I���̳�U�0�w�<'���8Y��}&�v�k�7�&����'�E��$n��0%�:UG�)�����ϼ$˫K��@Sq-f�ju�ff����
�h��u�����(�%к=qΓv1�� ���x�\>��C�w)���ގ��";KX7ޯ!Ӊ�c�dAO�@O���D`q4�$�h�M�g�h�O�R`�Tɾ���"1
�������<���l����{��&�1�=A�����)��浦i�䪤���dZm�ƀ�:����l.]}d
e+q���5lf�Rﭸb���|�|�ĳֱL�p
}8U�U�enXn��C�Pߦ�1��yR��b�{�:�[�/]@�/�N�0H�a@��g��ܚ-Rk2_uw8�@|{��(8�ͻ~�^?���Q�QOدѼ�ř�	�JՁP�yt��ٽ:>	5����B��s�ݸ�;*�q�3i��DO˘�_-��yN�_|�<Uj$aJ���4�{1�\׃���>�X�׈il��U||#"�2�87��j���Fc�n�$�U��T{>���;ሜ"u,��;2�B�ۆ�l���)_�{j�y�^&���п�})��K�4��	IЂ���a��~C;�\�2�H#�qt;��΅w�Z�E<'c,�̢��&l֒{�� ?y޷���Eq~�"��*w�z��/�*�\�2�p�2��#W������݉�����@���.Q����#1j)Rr�A`����&�8��7�yd�RhR����6�4K�V��$�