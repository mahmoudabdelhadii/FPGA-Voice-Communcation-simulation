��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���/�����Cc��<Nb��.�x{�>��0����=�����=8RLG�h+OLزV����ݗ�@��&�K��4cbXu�6@A��?��I�=��O�s=���
�S�i\��D���d3�q	��9/�I�w`W?ދ�S"K7��5�,l��C���
@E=D��!
����荾Z�V�h��c,Dt��&�����]4w9K_9O�=l�uE�w����[R�\�zÚ�-J�$����åCj�[�
����T=���K���h�����,������#�z~��?�G���B�~֨1)��k��yq�$/ju�YA9��SX�{@��mWt������w�F��r���������O)�mC�&�����$��^_��|�����=������A���_"�s���50��-�ݡ��kVE~�cu��'Ah%�����v2ݲK:|�g���7/��=Q�u�~��qC���
qSa�a�n�m(�]�h-�FK�]�Z<��K�b�s��'�����C$Yכֿ��h|�[@lXJ�*Qm?�аR��(�v�vlr�j)ڦ��0p�s�bv��jy�-����(��N�vהS��Y�n)!��\|9��;#�o:�#��9|TWL��L2=�'���$ƫ���19�?�:H�A���T秧���,rJ$�p}�a�ڡ�rn#9���~�1e�[e���!������{�T�7���O�z�������쉎�<o�j��D�7��lS�ƃ���F�V�:¦?�,�:4I~P�o6����2
�ԫ�#��G롔�qH���'> x������>I�nN1.�yφ�V�ǹW�)��	�3���k��c�Rw�buRA�8����\��L+p�q���ឿ��C,��_��6v����VN��t�["킐c�F�%^4�?�Z+��B�ϊ����o�
���������8��6�G��0�:���w��$�2ßt��q������ ����]����㜖@Th���oB�O�\���򨚋*5�2[�[8�$X`LE[�~����&��4��؋������>W�v֭��iI�ںL-��@� ������e^慸b#��]�Ԭ�|v|D�,om�@�Hr�`�bb�z 숂`��@.^�Z�)���F�|ƽҽ\�u�K�k�w~�%�/y��m�ً;zp:�`ʛ���3W)Q����s��b��&B��~��u�f�j%A:i�0Z���i�	�k�R��R����m�)���\��7F���b�!j�����^~?�!��G�K��#z�j���{�jZ���V�n����B4Xw�0�?#�� \��Jg��)���){�^v�nX���dQ�F�/�p�q�a����g��C�e�z�!���X�+H�]a�py5��i!�.-C���(�e����T4 �p�Qj�������^��tv�,��I�3�ιz��e1#���7�6���gY��<��d�$�3�'b��G�F�x��K��NdN/���"�b~�"_쯍[��ۑ��q����QB�A<�T4�ƿ$�`3�3f�'f�z���Y��<{��m����mH�0	`s!��r�ʴz�M�V0�AqՇ�P?����RF��eWH�=�ި��~�<��H[� ��T˪�k;؞R��*�p�'!`K]�;��,B���$H���MƁ�����*��������k���嶗Tmq�{�.H6��x��A�U�-d����H뭄a���ΒF��t�ϳ=������x���3Г����ĸH9���z�~�H�<�U{�J�A�Q%���O�� ��W�B
�Q�����ڝų֭g��Zj��ICF�cO��[ѣ�$�ixS�._J�T�Ē�a��I����$c���z�~_�+i�m�PW��6�xY#����t� j�$V��YoI�ۘv���d���?\�F�m8ǒq�[!��	�#���_�h�G �����=6��8(���ѝ� c-#5�7�̵��i�����7pb���2����S�݊g}�3��U�Tp7Σ�Pкm��L�|�ǸG��O=uެ�.)����?��`ߎV�H>�>?ܦ�0�c��4H�ŵ�-����i�$g:ڝ�2��]��i�a��+&	P��v\��v�d�a=�ۻE�����K��S��QS�Ǩ��@��X���X`�U��M�Z�DYo��a2PR���h'��x1wiDlŅћ�F�f���1�$������M�g��%y"E�C�Ӻ��A
��Df��]O��*N;h�AI×�4_NEO��P�O?��9ZB�̲C���\ޓ��X�D2m}=ԃl-L�����U��W�
[�'6��=�:A��_`�<5����<�u%txE?���z��w9��a:�.�!��2d7�L�=3I ���։y�c�3��k�*�����1����?^���3E)�w�;�Q�����1*M��H� �/#ƀ|�SF�t�X�i�#����*/
PGQh��ף��m�<��ݰkI]}���a"��C���$�p�4�����}>��L$��.��"���E�� ��#�#?fT�;4+6�=��y+�$��5���cL�)Y&�6��tb����78M8Q'����)���et�03����������HÆK�ڛ`�.���;_�����f�����<@M�*�=�O*�I욗j]LJl���Xˋ�sJ�3[$%A��?OD-�3f=oe}���x3�P���������d�z3r2�K�g��{<)f��-&�oR�3������^C�S͔��PE��p���C�*�o�ё�,�O�z�S1:y��+��L'~�y��h��۵Z�ԎS1Y>\�"�
Y�7V�-�͔w�I�����?ޙt�̾�)8���,1��h�t���y��͍P]�N5#�����5�z}�&�^�51��J��K�b��n�򼌢�Qd��p{���_`�8���0t���3����)~&�;� ���D�_�$��~��y�[Qc���f���[��+`�G埻aY���'18�����sb�ɷ(�Mq*�<�w׷j�@ �K��,���,h�y��L,���ƋX�Z�#���p.��.�4��@F۸��k�)�g������8�82�t�,؂M���0��N(N����P�\�ȓ�p��q'�E�rsFOd���x�u����J ����6��dq�ì}����#j���7����� #�=!�F�C��,�'�7�!���&����m��bU\%�P)T査d�nZ���H�.�Ź��{ɥ/�Я��o�H�V��A/��q�c����r������������n�ػ��k��zK�r�Ӊ��OT-��&o)?k�$��5%WNl�mS��ϒ��SuU/���&ϵ��˿��0��BP� ���?��C����,BG�'�V��
��7�X`�w�Zd&p}����S�lB�ks��W��UV[��iY���R�\Ec�e��z�CC<���Vg��L��5�!��0͏?!!�;��v�b�oн팂���Z�W\�)4�F�7F3�o)�X�K)
*ɺ�v�gx��Hr�a�?����!�>W��[�I�`��!*j�|`�֧�u��?��/�kZ.����8��$��{L�h�� ���;�sL t�DxId�&��n&҄m܅{_;C��Ί,^k�؛�f�p�7�ߞ����C7�);�EP�[���ԓ�S�U�U�dބ�-p�����AM9�J)��ns>�����r�����9���5�&x�x�}�#�]L/Y�&4�Y��R��E[�C�T֨�P|����K��m�=����&;U�O�-��_B��;�M��jx� �˂����v���G`��]��4�����n�!��\����Z������=����B�wo*n6
��L@���	�J��(=A��(�(�x+~/a��L�9^��w¨w�Bໃ<��#��ˆs�T],H�u�;����}���gF`�1�l��s�X!%�^)D��H�����{裡 G�X��m��1���fec��[�֡/wK�R~�T�P��{�ʢ�(j��	�De2*�=?��a�LU=b�!."[!]�Ч���>�}� �lt�'����?�k����ɃA
�Nԃl��u��Ƚ����u'DG�,��U�õc&A�� '����难��\JPɢ���9H�	TuT,
��2�_G��| ��1��9rh\A���j��w׳�>�+�:�K�W��X���ƪA����ѐD�Ջ�߅5/��ܳ�|�������u��,'I.��ߖ=�qΌ����M+��%ʠUZuS�=�g�s�M�&>��g���槁Y���a$`A�&�xf�E"�)e��֌�ˋo�i�ͪ��-��j+����@��4f��]e��"0R�"�e���T1%F'6�^F[�ʱ�Ǳ�Lm�d����n��i.��xu�5mjN�+������R6�5�������N�Ȍ�����v.�)��E�Cי��w�l�ZS����T��~n��Ye2�0��O��5�8�.�|���	�2�b�m�楩<E>�ZZ�
3\k�1�a��v)>yiVd�X^�6�b�Y���շL��^s����?)1P@�;3���Vx�0L�b��vY9�k`��E��*�� z�>�^���[ɂc�,2i�1�C�����j��qIۻ�5���T�[����6#W�Y�CtP\��b9���l(�θ���3�����MS]1�%*��\]׾a����i�O��7��Nz�tMS�m��e����f�~ ��X�j�nۖ�Z`��,�ע�:���nb`S�Z�C�H�R����B�0J4�$�i<+�%o��=�$]H+£����ὡw��4��~�C��(|���[g���j���u7=�T<M-�3@��"M)P�.����G�xX�Zz+9E� 3���2�@���լA�{y�AW	Qٯ��4�aZ�g7W�{O��s��=�W刲t������j#hg%�~�$�ט�X�՛�u"5�{�ER�e"�â�e�����;k��u`f<M��T-��У�����%�]�A /���*���Z�ͮ���,vtk�)^O���D�.��o"��Q�̴�	Kb���� ����b�8�fU�X����/|8���Yd���2v���B�D}����gF�B/sQn{�˩���������&C~w�A��Xbo���V�+j�`:��>+<����u8X��O�T�2�J�yF"�[����h�b��bD���@��?�8 V&I�8׾�^?;@|X�P�XK#/�f'�
��S��LEYW��7%�ʁ�$V:ѦN���xY�G�Y[pXAd�a�X��M�@����D�i��t~]*�%ӥ��^]�Z�� �SF�#:�;�-p�@)v<䒠6�i��M1���n@�`��^/9%&�.;<���R���Z�0WK^HjZ0�;����|�ポ��(�D�x(�������z�M�^��M��ڃ��@�dH�I>{��C?�\�Y���<��y��b�oF׺�)��[��:c��x]p>�!��ۛª���@�Z�%5�	�mŶo5������p�1͂=>:R=���cǢ7�A�h_��^��Z�I��r��4�/�@�A��Z/9�5��&^I]����[`��E[nu�Ȗ�&�������
 �Ba��VR�����㑔��P,g�����q[S��̟�����q�9SGR�ٯ����;ľ�������o���r`�
�������Z6������>�� U#��":i����_��z������E�{ILkΎ(~m�;9�[�-���(ăǧt�飰(߄i9{�)��7�bd�
Q�(6'��
���t!1�ҏ"����+S=�D%~yʽ���F���CB�,��b�j{
D�[i�}�g˵lX���f{S)�eS<��o�V[�\NW�)c\��庼6�W,;g���l1E��U|�(������(l-��^j�}!�6�����'Z	ډW��}�����ߣ@�r�ȼoN��[�\.xc!F��9�]^5����*�ns�S�޲7�?>d�fB�޶SI�j��a�	�ʶ��_tb~V��kӂ�#1!ĺ�F�����c��S@xJu�\9V�Yn���4Bq{���I���5a�6F�+%����E�T���	�M,f�Lk���56��c7��l���h��n������i���tv�ʖ���o���z��Ӝj%��ʧ_tV�=:����V�0 ��U ��K�
:��C-2?�d ���2U�.;��e���z�R�s=u��?p�먤�֔��P���:����A�^�<�T��������E�GсTvlB��)f+��H��&`Y����8��0�
3�ncw�U�3���V.VZ~��ǝ�+I���f~�a;�{13�$��|�o,���:�);�Y��I#Fz��S�lI.����4��'�!��$_��rL��
��sC�^Ť���fEֻ�<�8��̜V�f+�1:	)����⁹5��!~;��P#��@���|�~vj'�S�9aN�[�eE� ٓ +�N��;/`���F&�Ā6���͹��+���1�E;�=�bۊD�'�4?K��М�cf�����)�N��\=I�G֋4������۸�^����g(���U��K�d˲����`˗����钠��s	�\���fuJM��Q���q��Ck�ױ�{�&�Ho_�TG9�����L*�`4m'Y#���yÈ�x�&Aw�q�K��R��ɱ�߃�;�A�
�虭$�
Y����a�C�z}�����ῳX�iwm�����U�Mj��.�\[�ހS��:%��6I�XR�/�A��_Bj8gXq�u�ŁYr`=%�K�����9�Bz1c�G�]f=�#k'���T8^���Y��J���K�ʶL�:b����c�S0�A{�����yD��b0^��@�Q���H=�|h��ѷ��6�m��;��u2�N����P�s�j��5rn	�/8�v�o��O�!�]9e���Ii�u��ć3�T���_S4�M�ԾE�����ϟ��ْu�r��S��]$19UN�K�+_H+�,���v,}�o���(h��p�R�4��L���W�M�sA<�Y���(d�=�L�;��h,?�@j�b^�E�煗���*��i�E?�;�B�P�V��������ce�qİ��Ї����S��G�R�p��GJ�m��w�ʬ��}��-��
)r����~�7C��`�M��ReDI+9=��ᰚƽ%�0~q��o�z�Kk&"��E�3Ņo�˅�7�\��6��"WΚ;�	��<0?��쌰��������ʫo�K�R����(�>��c`:}{<g=>�m̶�i�٦���눹��J]�L��<"J
-����.-`m�
d��dj@�os:屌�¦&]�#��s��o�--���C�Yގ��җ�kǓ�E��6������}��bb��X�ܪ� ����N�$:�	�<q�м�(�X�����$ͥq�5q��Z~v�6g�"��ڃ��m�kC��g"1>�䆷O�B�?�,DZ���,y4|�l��|s� a�k��:���0ڵ7�d�v������
ԗ%��=ٌI��BW�d�a砎���5��a���Ķm9@{zyns��Yl������L���:�Q�H�L#AZ�z�ҿ��φg/����"8+����+�UY��
rz;w�E�m}=�����}�2�A���ndI�"�cҋ����cGJ���,`W>���>:�
���Rk2ʹ�|�R�x@�\�����d������Y������X}(��e����蜶h��Dc�ם���u����1!������l�(�҃gE����2�NaO����kȶ��N��PI@־��W>j��EQ�2����[�ZA�#Oh�Q�-N� ~4�?�ǒ���Ο������t�<Ag�RH�}�B}@V*�R7f��W�=� �E(�R�xV&T�}��1�oC}�i��t�?>�B�{g��g���(��3V�$��x9�����w��Lu�{��A(�rv�A�#�����zVK�
�y5��������Ky��~d�3�i+W��H��w�ʢ_-���\ɭK]�Y�~ce�&Q4D=q*�W@��b�^��b5����_��
�)!���[�-ժj�&R��|+Ġ�ȧf�����6+��N|�ǌ|E�Y�������i�x��Q�P(tR��J�V�E4L�@�-=��Al=�|��b�R���r�B&͕�
����!�1�U	_=�Y��������ڏF��d�#�!K�Ĕ���w���jM��]��B.�N��M�)�[P_�
�����������t�һQ�u>�,���ta���g��������3ذ��A�Oѻo,ũ���(�w,�r�7�~:�=w��ׂB(";�Q��eUھAP��C�)��b��q|��9[R���7Es�3��5x��2��A�0#����#�䶲����