// Copyright (C) 2016 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1
// ALTERA_TIMESTAMP:Tue Oct 25 01:51:03 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
YxKonzBXktk05tPYhhECjKE4Q0IRHDsWNl61gyMasx9u8YWeLjL3fGri6cCJxwXH
8hJvflSEFTatwcsUJ4z6yz8OfjPUMmbSrR8zlmRwXtHNV684tgN1oi6yg5XLvsto
K7XTTQ3HEwu0KXLPQdldzQyH8H2xww8KnKeFVKA4qsc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7952)
auf6GZ37eQgKyxgTCEhp1bAyx9oA3g24gXs03YVtw0xdA3i+YosONlrk+Uq+6K2R
uZgzZTTtkDKIkHlsdjrqYUiNv6Tr80c9Uiwj7OAA4EHN6ntgKNmAtrSOrM/Pc4su
ZgVOaJku3oxVFD6Ol/poTt6Z7Ft8FdDH/7/Dn60QuNp8qwNw6GSIY9Nz7gGvfdXi
vj3Xri55C6irllKTEOhqXbXu4Lc3wLeNs5M3hExRwtLlbkR6hrL8Z9gM9ZdRU0yh
WjWjSLXsd5TP8WeRgDJNtH/Z+DbCX/+73yvcjUdNSKH2ANGoxfuqDyCeJB2bqJsR
saqhcO4FBLNyj681J1WyLFFDj7vw7m8z75a1CJA/49XMy9ysv0EVDvgEHplk9e0g
nPA97Q4hWVTIPl/QCRvoy0KGi4Z2sX50vAhhw1FPJUuJpJLIPljFV5yv0phOwB/z
ohI+i4moAFILlG3YBGKeE024TNeaQPid3ufWn9s5TC9uKZdJ6WGSspUXXFoezrjQ
XidfArvcL7uDxvsGec/hbaOx45yPUVly80LkHjXlxq9qeCxLdjkckDpF+3RU0oJt
VCA+tASuzJHSYDJ9fR+qbNxlqEF6cnHvH6kQDp4jUoIGAYWN4JvTutk20pQlKMeg
WcknbSsRWUaJLkPj/isFfoJpAuCuHNloga+Itluu5cDJyibDgck0ZX9jQLX7le0G
WY4L/MMoZAQaxoelkgorGnIr0ACGlAtJHYB5G5g5F32MDTw14w3WFvlBm78ufzg5
dA4rEOjlqrzxThZ4ZBWZgLMKz5fRVQhzUdn/8O2bejfsiU4pw+mvbia2aMT6g8Mr
avkDpHy4tmB2Mhj+GNpLhMYS/OrkcQi5+DUTIdsbeHANpTjgWZfDwo4AoPYjKB6E
mnby/X9EQD+xqfXj4Nasc51XfAiy45B4ygZwoxEKCPO8PTq21T+Dj1BTilPhM+QZ
a9a0GabNm27is0927/MOaOCkMmn4pxqKxvIB3XfhJodXOU6FBj10sySOvz0ZWhHs
+DWMuh03L1K4WupWmPadzpGxSn6/tt5FJLkXrvpulAjP6CeG43xgQo18qwSGH9ay
AGpXxkb5lcyRr3ePF8HXF1N7eJj8IAgVDy3KGX2J1p5fHt6f3x/nME/q7bqHGrGH
5C5FuX0TKSnvOGkrIKAPXO4A8in627hmqBQMUX2KWs3vNbBeh5Vy+onlruxCF1cX
gl3jX1ZzaTOOHn8FBOdyJQFgFk0FrfxD7LEzs8+9PIYzAnCe6Pw9d9QUrKlBI0br
rC4A3AzQI4gUQ/Nmd02Fb5BByHCvQskV2PQwbtLSwrV9U8fJzrzeAgIOdUfJndrM
juH3qoAK/H5EgBtIjVFK4RLky9mtbztv9GpXq+JikPQVsjdyM60lWFXgWyZr/7mu
1okMAsZIUQIyOU857UR3BR7CgCHCZqmVuy1f064MVdGJ69KqySe3WQ/AsdFPn4Zi
3Sat8W1kAPAFNJgEynhsD7BNdwmbMfeUzPRhKZ0Ao3VfYYdgtJjFWh4he7fm9krU
OnJPzOvVhLaQOTCSSvcBWihSZZc/lUlrXEfTaLR1A4dQS91NKEbNEEiJVfrr1sSl
hjnZBMaaSOZdUqPtjogbGQJAi+9KflHgCH3CM10G1GWIhdfznJf7cCaJTtg6PsUy
2WLcSkLY0I1SfKW8hCBL9PIh8HFX8gpKXF3vM2fXJW4Ie8xLkPiN06txONz8KQ0V
0SOKzH0tjWAI/aAJ0OH3yvf0Rsc5JrkvAFZINEPe2H7qwU7aWnXA788rsZivjAx7
Wz+zwvFCLK2nNrVqCfF/N/Ho2fLPJf1n2SIFHA1GeJs3UtdohUsss1n49K7+DfbY
ZOMDljyeYdzsy2otiK8QZC2hqEwdElka3BwLL0xjYjmKrsnl2TWCuSJpa2j/3LHU
wLoNGZhdFEBp4o7NNfQMWXsZzFP282KYtoeCaJUtvkDEwh8Dk690XVbY54sG+5J1
vW78AGL/2OeP93dnThHhBLT2NOXRVtdu6r2lynb5yU1fxx+yiv+gG3StPiLPLHK4
gTcUvyqrnbNL059eBsEcOEeiksC5sI8T9lVV0SjeBkRvFztNcvt209OLp0AyWX/8
G66H5QoXgRE0ErMslVtw/uKn07zWASu15EvynLBq35OO2xilj49R8fTnca7ugUrK
Vz3s0mAR7kOoSgxp+5LfzAT81B4rJMSayHm2HrIXM7lB35L8RZ2KaVX19537I+IQ
qaXt74Kg1hORlRV4Bb1wn29cQkL44G1dXmmaaWMf+P8x6qhRgr2koHiw9RAaYbwO
uslA4Igo3+NmxtAOrVZlTKXCPWKCUQTkMUKyb/J8cqy6h4Ur2BzF5U2YwZY00Ppk
EnyDLn5xZD/e0bwf2Mb+mPdKMEHKspLVJaVfjMFeYKdMdW2yL2n02tyYwN0hoNC4
IXOnnjYB5cRTNDQjH1Ri6wTZFtM7YOfjj1/BZadRkGVSUKdELF1u+2hIspFnf4Pm
UV01BzMHOS1DhDrYi2Ebvy+S2XWjNEAJb0HJBD+Ht7o99cemERt8+ONNed+pb9CB
lHeaUVzgyrRhHxaSIeRSd64PB7ancurCjlJwrPlf4gtXfkFruWYXzsymO9YSBBCy
rP0DaCfykM6aka152PA/QEmZYDi+IKG4cA5k6f7chS2wpx8+BlZoWW/Pe2XXDBZL
eXO5MomI+Gn+xQky0PbYHxsGZ9NyVnCNGv3zIuOvrLtQ14vcxUy/cM+hpGkCYRPY
JMLBoNgc9WIEMwC2LcOaI7ZJIFMv5RxzjK1OGuTuNgyqgEtGkruyi33SSVDQIWA5
ReYHGtVxBmjMj2QIsYQJGgReoJwEg/OC0pAj/JUQqgN7OaxG4AdxQQZowGKAZJl/
sub+DOWr+wm5vWAjQoNhbUzZdzeAFcRYq5LVXdXkrpcTZZuZZYJvf0fB3CJhMPup
mm7bzjLwCf+7PKTpdki9ZcFcBgOXIVcrSIurFVTb6wYRd+bpF+EuYOR1EmAeLLkc
z4w1rAt6I64+QDGZyfLzpoRveWEu7MoRDeiIz9/xoSMsp+P2IesCiBvIPXK5RXuR
+xpZlKWJhjeB19Q6/h5hlqnJ3O480GtmNGmN0f7oLgTcjHnvzemck1vkp3/DfMoR
y2nW8W2x4EhRNJmmcZYzMJ4FlkAf2HDKMDF1L0lndenioSUnNhQztCKr1YcfqYh8
Sik53yxunEng0a3+5beYann//B3siDkpV3VnwXjZu44wLp4rlgaXdYuJmmOuKYaJ
/8uT4Vpc3d383unKyh8tv9VHjUTkZ9kW5+Bf+OafhwfrLc5PywI68yC4OZ+bPPis
p28XeZZafEmeVlUI3PJl0euHexXHztVaszpsMIYpwBC4hxD5shbJr2RWhhvrO7Gs
kzK0pxj6az2py4zwBOwFGDj68EgE2Ztc5/nSGClCrpGTORe7rKZShXZ7DD1swuMa
Al7AiZ444xc9DCQAhDcTGBDSYHez8g4GCj8qWm7cKq4RtiGSYqnOB37mlq9bmWfT
3rA1OAqjmHit7iw8k/QSK0ReQh2IZhCpw2Sig5zQ/sLt/y/kj3vfgLw1zxYYxTrL
Xvyzqz+9bP3F0ufFMbqMnsHOr5GmRScYdU+jWcp4tUJ25aHo2C9Lj/tXF645cv9F
+5W0epFyjfn6GkkfAWJCSPog9xw15N+V81h31iUlzWldMP79gGfPPdAjYXXVbb+m
91qc0J7okh59k4ss6wNtZPkmsdmu3BV4fSrl9zAndhr3mlS2LtCrQULx4Cz1DMhz
pn+qNTx0Zcz5tOc5giNe/E6zZknnijMnk5lz5AI1rBoLwhRzig+RYV5AdE5RQuXN
PURbQu1EnURJsB4gt9Cz/KrsC6tChR82Wdgs7CeNWMqBAmI1KMvyjAox73xqRbOU
j0PWZ1yf3xns21kNjERnI33GQDn8vuUWZvVoGFt01IJ/zMP9Ha9Oa2XvTpuCofAB
gYjNfTPRT4c72Ywgo/Mc8/B9BEheAE+e1O2tp1WOJLc1l4ALXa+3NjvrJKDlUJTE
7IOJOAhwI77ravwDgZrncLuy5Oq5A8NJkRhg0gkYa42IkrPgkM8R+IIUePD7wdnP
dvFfN/5BhT5IWt/TEVlZk6O0BGIwR8GqOIf8IeWrSZZjCF3g5S0iuaV2CtSz46S1
rrEGBp4EUqyyvTN/F7i5AHadyXvqUlZtL+s9DQCIqGj7tobgeIiWT0h1lgP95UtK
92Dqvxh+UusS5T8eDQ25SihlDR5mQojCbJP994INP5WICT4uZLt+Pq43IdaAlQTQ
hBj87QRs/7eR6PjnmFnwMZ7UKQF7GjP3v/5G9BR4vxPAJQKKp10APNbpQvTMfhxG
z+RI8DFH48WkOn+cqEw6Usp0XRvVlnn1K/lMsJ6ENoNho8qAmaRCc6997l0c0BMc
0A9RUofRgvZ0tI5qMN6hu5ba+ptdssjjJggjNAaGgw8RdgDdswl7KADCLb63LP9h
PS/tEQ5NUuw13nUGPs2TIzS4YQaSsDImRyZvZBhc7gM6TtBRnkYKb5JfNo9CXXVI
bVbsUSn0+OWwzDgYSCve9GII2XSs3nHaqandqFg+KIhE2E4bmE4TFbjBl26hLmxp
qUQu7Vb2qdHO+C0zj1A9LrsasAsqG0wYp7sV8Tepcoxzo0v+2Kmb3KQhx/2fByok
X/bPjkAN/kihzLqiu+vwzt2sbveikHBhrrmih0ewmNnMG9jOtlfQk5dVHZbIUwEv
h99ZwOtRubeWeqnRF5g4Ojd8m07k1YgcR4IuJZGHIpb6AJecPHlByvNcWcJBMQ15
W0e19yOM103flwTKPon0Ml0aTn4rGwz5NwN7T0vWtC1BCOaAGiDtGo7FKEzx9pCV
Ed7QNbADQMlTuq2zY1TipMEExmFceYt5Hrv2tINpMuJxUjjifkRvYijT3iJtQLTz
GK7Ti74FQwrqYUxlwuY8kuSg4bnzPlOW+Z69LVV5XuJWx1McEt2F/0efaqXGhAmN
u3iQsyiH8vKRE5ZbD9evoMAjKaV1uQnZTZmqRqzD7n/P+yRM6a+4GU2Em2Yzrzp1
QAfPXfBokAtrOvxuIWj0eDpTcgYIgzqe6YzkZW/t6IjqS7quaHerhul/bytxIGvA
j6Cyb/T+EwZjlit680ic/qegTuDOhNet00p4UEEX5N07i4xKac83Cw75RyzFMGFi
M9LidUNMP7qg8vxwNLoHxAQ68ZBXrLyflSUCPZ11JxkrOxHjv2B2ZWoaDyvahF36
GBs+Zo99qld01cD6UkqD2wSHT+mBLFN9R9vHoexxCM3zcm+xaLpSqgV20bQZmRMD
iXWYWAtSGXNi438HlLDaL8q6R/jFjtvLZDoTJKQNefrfOsWbDrp2rDzCRzMH+f27
NSF30bjmgiH+plKtED5q3aZmSYDyjPKPdWm/65Jrvqe9FUtN7sQo1ZUPUE+9aGVQ
girfx7vFcs07wohnA7uh8ntzCoHfzSc3Y5KZ7QijxuTxJ5EM21kvcZqJK6sIM0G5
yrPJDOMcSS24DecDAnq2T2IDZDy2qifp75rTMfqAUVey3Fhx2xh7Wn8+vBZDPwtv
061pC0cDxQiojRSM3D6poHM5TXTtsmE1Sh4UTtTkxn12ZQ25PvkXg3A6zdEuvm9C
3QErcWNxSFdRAF/AG92CWlECFovIpRz1DyQ/i6bwvvSm/14xIc/i+nBicdCTxG0R
wX8BjHC16PK5LokQPO0c3xB6nVxsSIojY+P4JZfwLzJZwDAxJJxZFAwOLJSnDSZt
VgoJL0Sr9B+ZpXdOQiSeBR9erghVEzbjCFJi0UmJmkaMxW1/IBFExZnswTmSYsND
P3Iz8TzGct7q43UCkwgAEWpwN/2F/yNoXYS90obYCElK+SBK0CKxKDR9vSCiBupC
GT6vplGs4ynBTwPuRobT8ViLuNlnLGbDFfcfwo5tlcAw78dq19PtGvdiMZVsowVb
i9gVOHr5tRQWtSy6hv7Dc3qfUwfSLExAzNqR49lGVFncBuZCiNz1DeH821Yxs6dz
bFO42oV33amGu+YdPxq02CD28DIj9wELifoJOeNFuYdgi+6hKw9dkZcTDBafLwok
VdOqH2sbgfIbiy47lgxF0T9c2IebGENhcjqguqRfLmf4/wVkLlU+aROIcgCSQWMo
5RtjWeof0KOIvAo3XXT+1nI5pl7RWS60KV6inbSzGYjews59yjMesFXhS8JvFsHn
jkGUmYImTo6WQYdcwcOcr0ZGqXo75dDU2moTXV+/FdNKsdvMml6mFHNoNPQoX3TR
NbVcpICJ6X8t3OMTzI6QSuwUjEBjwvfFpxGd056OfvozQtX4c3WUpUcH1v3BHqk5
R7b1MWmVlI69i3p+N/qX1IQKv8V29AroSlf2vYS1D95U2ishp6LGD2vBOsnuSItx
wBYm111sYobr44xJihf4+42+A8dQoBcCMIH0yuuSz6Rk7Mog9U/UqB3clnHhgXJp
HUZkyKxw3qIJ6z14HXC4g7tZMHwfBSTAO76Anu6T7LuRWP4pfP0hWQB3U7ydTKuH
jDA08HBQ+Jk7t+x9ohlfexrZ2kaciPI8D6WJcDHXIXG5sNeGs3/UDkh+1sgbPglR
yXnZxHPrCCKta7edB5aMuWTszcJV13c2NC65f0J95XG1/Dpf/yiVSiTUnotEX1Nn
fouXdxlqCSsA0kfWAw/CuLU4ctxIlgXt9gNvciz1TT+fY+/I9ZzomMm5mIzllYk8
aUKDlgBFG9hB2Iwq0HeTnWwM5x1SFK3yP1nyG39gN33LXnA7OSCjxGVVaYrLITXU
lZhKhIYb5voXkykQu47ZzskzRZBA7otnSIvXbmI5ZGJtH40xmC64Idag4ec25smz
LY1zcfrnvzjKe6XnP5mkb6od32L3qu7eXpbPUMMgsGA8cIoAs2hdongNh0mV094T
SMGayrhP6o+qKaooeDQk8C/SeGYwhyVSHM+kJshN9oAuW5pQjAOcQfcc8W5sKADF
2MdVZ1+2aQ3O3d8jZckrtI0Qo2KFe0FITX1knrjYrieG49YnlSDwaTnSxNQbICF+
TQpkDY7fKpU4kJo0pMGWwW/gRtjwhrMau6V6T6VOpMwTaz3oBqeaRNlPngE0MmmL
creoS+rHNt+9Sj0JFYtiF7gwROBXo15DCCVfnAZZWkW/jENMwL8qbppe9ciyPSVG
xYDTOqEX4aAhwCEebaCqCsJqxTxqyGyEiETdEKoxXF3lM/vBjfM6AwXk5JCz1i5p
ohzKOL0VovF/j6XNr1x3Yy81zUrF1WW6MlCAv6Hcy+375J61qYxVozW8825ZeBvL
OsVBW48usivO/dVQh3OHiHzLE2vhz5lOfNRm0CHrUDWj9YlM0Yb5dded2DYowq3n
7ksqjf0Ywvurb6WSrLptf9NiBDXTFlm5Od8pzWvtczg543JPUn7K1osWWi9Ytb6X
Py88QNdVlFW2xd8erJvff26Z4gUFUNYzq8Eyu6XxuRjWJEqGllhZ5itlKW71c9xy
Y0S16Lt/jVMcpUe5yR8fbw0bEceVOK+w8pnObh0euiZM33FskWUKckKDhEH8n4Gb
Odq2XRfBIak12TTD2M1UXvhc4/HpCPofZGmOMuKHAXZYwhNsECJSEoxXg6w7CTTq
n4biXE3zPa0mpgJUwSLAkmmZ7btd3cP6YsclRCYcedCnp5NwpAxdwVd5kKFbSb3J
kOCFqQwEWCHdh3i6C/6VYBPHeGzTn1aTMZz5cvCI8Gd22VA+w/5Eednlwlr+Qj3M
AByvhS+G/V0hHmNRDXchHzCaioGvMe2QcP1X2NskBgkwMgappeRbmaaPBJR99ggp
X8TinF5/4qcPXzFVy3O89Io6ligmU3Wzwm5hACmkUgUYmCpRbz1HkoksDILTca1N
UFQ+2jyvCzOSJYWqIDt5Eo6LsE6PSK9/C6KISxBa72USsA61yebiRTztOV2yiMHQ
pUtpmhvN8DL+rmnKhFIdQMGjGwwSz7WBwHEH9RKfJRluZExCJziTymZvlD9PlCt9
eE3E1VSQRxVES3iTMC7oR5aD6MWymMMiW1qzJTuHuObIwxAbaBGxTZK0QVXAzJxV
XdwDTzp5qbUm5SNy+Qzh4jrvD1UU8BYTGdes1as6X9+ughWRMmW5S3dPT2pCgPf5
nG/GH9VXoddGaO4e7ioiaigZGZOVYOOBA6VA5h0V5LLm5W3upqVH40HLIavMz/wd
xfUbj0F1wYq9rU7JH3uL2E9eneJ+2AeSDbln82fJNpghvQgHQqm/zB5lq6H6MCRr
QwFEBDxSx8Bmlv3+tw9R/au6RixJ5FM7vwzPlfAKMy4annyxJmbeRv7QM5bFgCJO
HpHyLLUCa2IelITyUq9YEiCmyYkb4uPv6KSpE4oCC2Xk16qmwj5cZxbRgPnf7qwU
Cv5Lq2iUNypYHtG8HgkVQJJ/Ch2Ne5HT6TT2r29bVkSbxHpTODNMDenYlHGgL9u0
BLs8Wt60ThMbVJ6PEqBTDU24SDZvYh80mrvytz8XeWOuaC21vwUQLhBJ4JQy5e5I
EiFn9a/m5M1tOflWYfjOUaeBN6MbT8kkCZnEzvkVsMOvSRDbfJqfjYHheOWFjeLo
x7xBMauLSExdUDvChRHi7CwtFFPt46oUx61UXjywI8zz6d4aQDS7dzNV06tdwIxk
g48jUysmGvdBi5vezVWutBnyIgOFXmbCCR4V271U410L0aOlUd80vLWBuLlRCuE6
ryLfbrlta0Lwe1f4yvnp9APpuxla0/R4zVYBdVx22MAvB7ZgZ9AjdOybBXdv8DNN
D7/p16nIDyOHe7VJ7k95zOEeqQYsyeR78kNQQxl2qlHvC6sMzlKi/8ZiE22DKXmC
Br/jT8y48nyiMBem6Uo0mqwJbadnG0d7tF3v5WvDY+ssFVXGqJh8aoV2BdTh8ehf
sj927N1Rl69olCFs9O8UcXgFKJaj7KMM24QoOePlXKv6LiskHKEzMTck86PGk51P
nW6qBSpwQPb4lr4rtoutfDsFa67I0X6O4nI3sRkVcptxRFSAN7RuT72jqAqYTPXz
NC3oC/dNHahyYSoI3IfJgAWDEN7LjRb1cN5p1kbQIJaTXcn5KCS3M+rCPm2wJxjw
27II3XMzBwIF1T875BbruQDTA97U2+QoG0FH6TeH2HdfGOWmUqRRL1Rvho2b3Ovh
7ibhBbfNz6Ceqt5037D3ZI6GAiBeYndGa+YjsQIU4sgH9yZOQl+fzQpzu9rjdBds
aHjGPWEn/Sebtumnfnh1iH9VgcmSws21jx/9HwhqPl2xdyeRb93pgATWo6gxt290
8HZaY1R4IBQSKd1NQcKk7uYo2i5RFG43EEVjiUrW0WjZGiH09XZs4P5TYETC/Jws
jxLfD8ppkq1oi/7cOSpUJ1V5tufaxwHlV8ZjEvwkDIlRBU59qmYycJxwln6lgYjU
bCDs+A7N9/kT9HJNGPOCJSJCC9yrwubKLBmOI2qM86Gq29dY7s5SZDcatheyyPMu
z+JV3Qyiif6xt7uHUGH3kHTr7vjUtfPWvB7WjBPBSqrMa5nJFLIjOcEl0ovkaQUa
VdJpiKi2czbKbc9hsZ6m0P2VHRezknq8Z2LLz7VNmqs6qGdax4eqsXy8bpnrgl8v
s6Py6loCnNFkjydnos9kesWRHn4MTKt5hX/hx4nZcMhzBpbJcO37iTo4zwE3zF54
a+xJ3MyXqdUETboiaKaj7zqDVeXUZNIo/m+wv/naOS+mCG9PzHSuFY1lEIpkvAcU
ZrGNURkc7qu2DbofNB5Mjfn3SmvGWSuVLlXOSn+KUjOhziNqyVwXWDAropdqRsMX
9gGJAYrR96k/T6PkH/7X6/8knEDWVoswSE6BBCi51/kW+NXahNo4A5h4+eL3yArD
jJQk+NvwwvGsWY/vg/N8X8CgSeU8QMH4B3BleqJ/KnpK8pUrf0rv3T2WT7bYdsvJ
dUZ0QQ3DQ/tmZ3fJwTJ+itkFWYglwSV5Y8bFPLAlvj/BLsvbAFYd9SJhvLEU5Pnf
6/wcAObsaW4xlTCAy6AiHEpFLHZ2+dDsGVFJs49qFDc9qfqpaZtlXyEIoYuNoahN
afQlyaiRYEr/0qnXHHOSwV9oMUV36XmfRKXCsxmQQsWdQBzgbmnGIIrIJ63R7VNc
FR/thnYHcsEYVF6hzrWDpYYo4XMYabvZoUdEd6QwaXUcyuCSX4QA7dg9op6kJRge
X8qQWCDhvPHRwmbmM6tMsRP5FxypCweJz0H8nWoSvb5pnJoOcTCPZK7Dh2XxefNW
uC7Z0Q5RGaOHK5cAhFJtBVw+rF5gRqrNFFfTSDrpFZ+GnY81Pp64lMHdr+niZuwB
Do2RGO8Ok6LnjrfpGCgvdzaueX3Fh4JzjbCdgzzkcShAUM0zt4g/r42EvKgqPfvo
zq16LU8agHxBH4t6Huk6ZSwTuk7otofBAaKxm2BsYhq/Ng9V+wuF1aRUqCaRP37Y
5I5G8ggKTZEu6PPj3qLMpn4nEq+Y1CtMQ/OcBMe8/Cbo6vTvXIVXx7CU/1cu1wS/
NzU9NN3fs/v39M/sE0+fbtd5Zj+NksV7e8+dAjOtp98qx5WktSh2UJNyqTUzsAJ1
8g4qLgmSDYv+qEHW0KH2C83PcEMi67VaWXE/KrgKkgE=
`pragma protect end_protected
