// RSencoder.v

// Generated using ACDS version 16.1 196

`timescale 1 ps / 1 ps
module RSencoder (
		input  wire        clk_clk,           //   clk.clk
		input  wire        in_startofpacket,  //    in.startofpacket
		input  wire        in_endofpacket,    //      .endofpacket
		input  wire        in_valid,          //      .valid
		output wire        in_ready,          //      .ready
		input  wire [79:0] in_data,           //      .data
		output wire        out_startofpacket, //   out.startofpacket
		output wire        out_endofpacket,   //      .endofpacket
		output wire        out_valid,         //      .valid
		output wire [79:0] out_data,          //      .data
		input  wire        reset_reset_n      // reset.reset_n
	);

	RSencoder_highspeed_rs_0 #(
		.CHANNEL        (1),
		.BITSPERSYMBOL  (8),
		.N              (255),
		.IRRPOL         (285),
		.PAR            (10),
		.BMSPEED        (4),
		.USERAM         (1),
		.USETRUEDUALRAM (1),
		.USEECCFORRAM   (0),
		.USE_BKP        (0),
		.USE_BYPASS     (0)
	) highspeed_rs_0 (
		.clk_clk           (clk_clk),           //   clk.clk
		.reset_reset_n     (reset_reset_n),     // reset.reset_n
		.in_startofpacket  (in_startofpacket),  //    in.startofpacket
		.in_endofpacket    (in_endofpacket),    //      .endofpacket
		.in_valid          (in_valid),          //      .valid
		.in_ready          (in_ready),          //      .ready
		.in_data           (in_data),           //      .data
		.out_startofpacket (out_startofpacket), //   out.startofpacket
		.out_endofpacket   (out_endofpacket),   //      .endofpacket
		.out_valid         (out_valid),         //      .valid
		.out_data          (out_data)           //      .data
	);

endmodule
