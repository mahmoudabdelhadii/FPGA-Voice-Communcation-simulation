��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��,�y�}�ǰ�=4d�H���`I"��W�`r���T:tB�T4D�m�)�	1��I�t��
��8(�8t>s)ו�."[�漆���]�~�]��;�O(1#5�-� 偙O��QZ��~rL'�x[�i,mׇp���O�I43��4d�,�H�����SN��d���3���r��m���̨T�I;uj2Y� Er�*p�Q$Gm���p�V�`�2^���,hz�<p��l�Bxt�5��s��\yq���#�@W���f:m��T�	,*�񞭋����_��㧋l�	�\�:��uGd��PǷ��N�I��_����Tuv� ���us�(H�~�{2H�:Zor�Q	#%�3ˠ!��iS��95�,?�.���/�F�i{#���Tp5����Ҥ0{%���2vpn���X�����@l����3dc�ק�3	�Ed&3�ZN O���z��s�yxӡt��v*}ԫy nj#��lc��m戭k[��5)�A#�����8�!�]�Z�s�M���t��w�!��'ÒE�rv��Ϝ�c@<U��\tq+��&|�&X1)C�����r�A~��B�&�����s�:n{p��͠R�X⺂L^��R����c���f��J^?��ܣR�O 1�rV���:��T�4���AD����˩�F�w��)Dm�O�b,�a���1$��c��7t[i2>�ޔ0,S���󧇳Ϟ�ᒨ�-��}�!6��Jyv�醊�^_�(�H�(y^����o#����X��3-�k\8�M�T�"`R�DF6ȕ� �,5�;Ҭ C�k���1\������k�t־9�}���� ���QHF��"��t�9 ?��{E_�7��!����](�S��0�q��w�9��=�i]�1�GʦȪc�W�XC�|�$��}q�6����zf(����լml�dz������*�eLD�*�,�m�]ہ6����D�Gw� �g��' A���FX��\өܹ&�6�h�Ð�$�(+��埧��= Eza ��찠pr[�c&��nP��x�2�TK�M�V���3Y4vIR\������ɭ�1՟?4�_y�y+����ƄJMm����@����m�����c�t�����:ud�Q�����T4���QxBŎ��\o���t�*Z�$�*7<�t~eP/`lfhg��6��[nn��#<����n�D:��-�C��t��J�.�^kʑ�L�2ّq��M����ڑ��0�O1l2=�_�tL�\�^��YB�ŝV�*��Fr�m-jb/R�T-+0K:����
@7&HB�b��P���u�I��u��TFq�uk	gv"(X �ҟiDz5����<�����k�P0\D�:'��SZ$�B�F��eu�N�z%�^�K��b���i��M���*�s��%�:��EV�^�3�����c�Äqmy�$�̣�<rr�R m��ݑקA��&]�x�_5r���a�3�ɒ�#" �G��jc�ůi���<�ns��]���wR;� 1�V��?������p���L#0���"��% ��񮑸F���5�����X^�`u\���Q�+ƪ�e�d=��V�oIg�h��q�
�TDEр|���"��������" ���-oZ�v�/�����;� �������wip�d�x
+�+*�9����5^�fcq,���1wH�����?w��V�2�%[�������Fx�(��E���d�]�����nq���Y�2x>=�>"���w��39D�%��0m�j��Z,�c���Җ��"�϶{%Զ���/�O�TAm�HصS�O�����pϦ|H̍�L>�$���U�S��r���,�plV�h1
�K��� �O�����ә��D-Le��4����*�A{��px� ���A�w���;ϔ�HT#��Z�~t1�t��"֭�߂�T�ނ��/+Ý5�{��H9�$���޻��Ѯ!���H����������o�bB��A�g��n:;�,��ɍ����!��z}��<�g+���r�P'TwX���U�a��3�>{^J<<T�$��.�7<eW�3��S�IWpIq��l�T���u�7ZTά��d��D��<OG��^�-�]zv�s�?QX�5破^Q�L��B��W��[�ߋ�= w�$0vׂ�0G���\��:^�W�������X���`�HPH�����'`���JL��N�Jy/�rI�h�#R�ڎQt�o��;���	|*��*Ѓ�����H���%a�?>r�e����Et=�۹�ǳ��7��(��+����X<�TFhf����<<8� )��N��s�3K�z8/�ME��L4���Ɖ�3Bj�w��_
Vv���x��Fb���� �oY�b���1߈!ʪ�w5�t���U8W��ٴ?��|���]k¦���<��&����q"��k���X�*��K��)�-��\�)S�_�^$�$��F�Sf��^NԶ��:�WQT�\�9��lB�t�����ip���sx����=�5��4�t>������a�m#Ќ�����w=s�i��|��c�����f�[
�@�1���Ԇ9��
�*$7-��_hJ�/���\n��<+�|��J9��Y֑����kT�sJC����p>�rff^��m�br�ˢ���yR�V�Z����q������]�
�N�����y����j������i?�hG%����6�i#>�!�X��#핚�Sl�<Q�9�2�S'	v���Rr�j��?M��ܮ�]�_�s$'��R/7��k������%ɱˀ3ҋ2I�sv���r���T*� ���됀,�M��)q,�_[�H���5h�'�`���#�۟$uUHy��YO*�r�׈�P@���e��@2YO�I;tV�j2���FL�cp���#�v7��!uɕ��?����;����݉U�#N][�7p�C�ucn?	�>�Zl�B������2~7o޽b�a��� -|�bo$�:�w
G��vza��]r��Y����]�Ȭ Ό��i�����"�RvK�Χ�~jI,-�(�\�(P�c��uu����=�1f��Ō�q�%�9V�h�}�ݤ牆6���q���a��M���
RX-e����-��ґep�E<Q$�c�,�R��q�
|�s�iq֪M���?��ź.��K/�����u��|�Ay�����c2p�D��M�������e~m徭T�U���!yh��˭7JR�ῃ�X����K�����'xw����p�ټ���UT�2��D�oAA���ZM�0�>��!1����^�wR�r��|��֒�Y�iSK����BΤB���S�D�Z���mK����MH;&e�ɬnL/BXpO=!���,�r0{�������N9'�`�v;$�&���Ɨ �5wqV ۶D�t��F��̽�Fps��QՍ�\zA*k�>�(�=�R),�`:�.pON2?Ӓg/8z&p�� �f�H,28�a�oi�3�I�	u�{�*�4X"x%8��'���O?�տqqA��+�cr�Ef�y���+� ���ω�B�������w������ h �.�bо�r���KpI��N���+��!��4e���}P~jQ�����A�)@��A� 罋(>fY�ç��8x�c��&&�)m1}5y�a��,��mߦ�j^����^;⒭�����W͓+	����;��f�i�L��S�����05
(Щa*�#n2�};�G%���