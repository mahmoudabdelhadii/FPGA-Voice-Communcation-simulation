-- (C) 2001-2016 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
gqq24oN6ohk7DUjE0fugj+m5G+8mxyfyP9XBke71oVsk10S/8ErcZ7JFTLivwKRvADW1Wg7U9LK4
rjkCUOGXlge+2630PWKh05wvgrvE4CXUBbnaOGUyP01gY0hc1M71jymFR5zRCUZ8L/Mc+KQvCR8z
e2Nwy5qzE8cMMRgMWf006lAcBwWZZNZf6IlG520EQA5Dsu5tq+yaUeuhBsfDLr5es5MC1RWBVtJ1
9k6XRyzEhUqw9Pleedv0W65nodT34SJjy+45VLQkgnxNX0jDzHwGF+q2doPvtPZBSaKuXqk5fKhe
YnsDjxa6XXUA9HoRRZEpE6OmfIbY0dBEqQTqjg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 8160)
`protect data_block
2DeUA/8bUAmOa7dWsAFppuMd8Y8afijDFZ0YvTMWab41huCwNgftjRBSlPqbmQmzWqSJLltGKFve
5bixDZ+JkBJZwb0EfOFI7p929I6Yt9WazuBDVzEtzCLOgZYcV16sWZJ1t6Dby1Cpf16VLGTGD9od
ieU4YU1/aKVzmZ8GJA+153Zp9SAbWu8nnNzGF34xrhdt2CyZhJaGgwMfJBs6VSwhoziz8PKEJ8gR
BKMvRW9C+RFgQXo0/fCze8VsbPiU/sbrY5E6qHqGxdLzpC0gz1sZpZoR7HTOMF6nDJLBJs+0DCXx
S9VcpQ2Q1uRAzacpyVuL+p842Ibjw50K6jBwk5nbvLCMl65VVV/p3Ynd9+YU4xXieR+KPR72cjaI
NCczsso5LO3qLpLBl9rw7nC2q9zZ/zbnkZoKIrslMqL0o0kl4w2z2dcpPKVfxFkkgPReWeysE81C
c4jcbSWNbKuyuqBuvE67hpfGvwbvY4lhwjrqPQAqpOBNaVjFFgH7kkf9m4QKjqd9rFXoZfEJX7Jp
8nZScP/5RKKiMIodZsZfTfOti810AmIWsiKrOo2cziUIW3rnpmOR+39JfQrneuHNRjywj8V63Dg8
IB8YyIFjEfyrPnCGOSegRoMz/IoIXOERAodZZ2xelg5ahdG04ac+GwEEXZu3fspk904WNF5wXWh5
CX2c12ue2n2ZgA/CwqBI6yDRY4UBV6/SivKJZPQpP1PgTr75in6fS1JvRy7KbBoIQCFozYwB+Nrm
3VAW+iV4Iw7QKcqiHcCUGFZI/HegGHFgCE7H9UOYRPmcsi8743PGqh2bjI1SYiR7bKp4CyD0MTaz
4FF78Rj9ipEDjYF5BxGff9VibBYj87Na4ii1vupaBErw6GUEu41hFOJjU+S6WZhogWPznNmT36mg
NFwM3hIm+9zaFItmz9LjYns4tgAN1z4WiDAPNI2F/BMYonTW4M+ouh1f++LHMGe7nbzB31zsp+Ns
KSe8pBT/D+FWPeSWpmCxUJyysxYgdbO2yhAl9qTpwELO5bw1/wtjXkUDc2kj+/SwfCOS2BHByEZ6
m6gQzpB8QNBg3a4kVnT2w2u/wKR86at3zVV6LxVmfhiq+HpH6+CGsP2GJHkNf9XPM2XEl/iOD0Xp
Qz5N8weOP0K2CCgYEWE+WKtAlifG9Pmhum98gaPzMU6eGeH7NWnkDiAU8FHeASMDlIoroRroS1Xv
L3NiQ5whF0riwIhkbW2qyCwwGc8Gx0K3N6Otrsdim8biUD7Q3lBWP4wk6BmLmrZI/Z5PwUVLiHY8
wTvuPmcbTUp2vT4V0rlvwkb1UGAIXTlIMyhnWK8FRg8M/0Ssic/yTL69rURHXfFgndiMqBbx/bua
lWt/dlONqrd2+lHA1MCDgfKrYOvkov6sYreKSR5CmAFtkAM7X7fkSWLkuRC9EYR7iPq2TGb6LLPG
OpbcE3Ihw6pOIu6RWn8vrRAJv45+HxbuOZYyEEgKOnGxeCvL47P4rPhxKQp0e3fVfniBTkGDHdV6
q9eZBPJ0TTarMG5Vy5D7bWn0MJiRN0AhPC3q3vw9hwY2Td7EGBJx9UvultOwAak4LGHbR+BylgBe
YVNsGwk/pRCM49hK8GYLVpvDM9/LDREw5P4Jzv9lPhgxKPoluyNglJyrBq2CWfktBAYzAPflULTY
Zg+O9vMJh3vlXI+3PhpLlrHVdd7hjHBEM3naoWUQ03ui6EEvErXu3tLHOlq1rUwKR63NLIpXiWdu
1f2zcyNnYepg7FrOqLA6Hnq2Bx7BoJmeSOMih9/P1w6b+sUAvdIouQ4ab2oBLXKp1ZK+W7X1biuz
7HhvysQ/ROVBGVmWp2PbC24YrtF51PxjOx9j058GfERWu8A+wVLMLgmeu6pyUX1AvsngL8Ld7Lul
Ln9z4aNxfux4OE4XjBTe/64aeLULfEexm0LdCG0VcoFpS+W3YsJl+LYpbMndVEvsgZokIlMbzMhI
WylkcBhRqkEm7qsY8as2dsHINJ2Bh+3S+i2lyLTsCX1vvGewNXkQt8G+8NSwj9xiHUhxmIeXRtS3
qtuk6AUZzigWq/Rqcj/13vNZ4D3sgd1bldaAHMrYhDwYlby18lioFWqbyF9IPgOyGDuKiNGkXW0F
KuaRbMqWsAA0Yul1kjjPxdod/fgmHPislXMCxUamhGgKEDxeavDOXPZA5+Ord7o+aX5+63kg7A6u
+8eQ4YCRkkwseLfXtNS0JpcRPRf4PQzMiY0Gwl4o96fvI3/PnCgTAtLKuta7na00rllPprV09oXm
CKto+nrMq68r6Gkz5qNBWaxBZXDnXReUWLKJie0KKQEM6YAeK255y+VlVVbdEhgsfq95558ur6GN
I780NiGHTrwLYRZEjydLRKKiH+rGYpRSHTPo5UBbTXTxm2fihkLw2QcRmf1phXaZHbyXS4Tznerb
5+zJIszbFV5BO8suO/lVvfCn8uLZfnsPQXxFzsNjajCqFtmalwhYg2jIIi/KLVFKpwcCbxlbplf3
m2sI5V2uqEXjefG9EU2h1+w0Lt134ZVMWXYeVVEcQ/mVpOzwccUtE9i5+/xQF4gyUq/uFQJXUXmd
Jv2n71Jg2hiZZv3l51+/fOA/N/Sdp58jhbAHZ43ExMn5Afxkx0lntC7Iv5PQFzOiv5SNouDzaN8X
I8DqoE7iZe20wyxipiLRUZtVRGPGPFBaABEA7HTTq0mHJYfwWj6I70WHwiOfAsIl44jtQplwzCSE
3qE4ju02X+wOxoOUjLEtHMq323MiQMG6x0L773+jVCoN1kodmrO0s7QjA96zUjhu45hmkeipgBcP
eXBFnNUHC5utb9RxGTUd5QWp9O15xBDS5dX3bCOkqN0XqIR6FWtx+Qmh0gZ+N7NHlGOyZIs4E2V2
mYzxLGKaXRI+gCmfZpllXgmm+WVad5Zyurs524Sdg7xa7mQsjze78+VUGDxp6aUzsbXb6guPkJKv
9sxJT30c8p+rOStD5tbeqhkOG258u3cbN8nkfP74ENPX7+fJMvn84JJQqYYrH7uB2DKxHez5m0yY
CUiPklzJsUbqGSQX9+OjzfQf+0/4TW/f6CQzk+MY4UT07ePjHELnX0MCMCDuG8NtCrFtpUZnrO7N
ilOt2R0ULeqYmOO82GHyzshpGT5SMxd/cyCxXyz2sDSC6F2Y/2nNKX79/5ZsLERUkYhSRxslEwpy
imjL69CoZsbJj/u4lsO5YWFM7OFhtS58oz1Hind7oNa4V7EfEw1DMFAFmakLQC/Kf/f22ilg4qBh
ImauYZmuISFz2SfCbbIwHcBCRnC/YqvmXSEQwCLeM83XZ9dTNOPOzL6PEEo84VbHftV8AOwViHOt
9gyUsmavwzgEzGxBHuS59MbRngTnF9yXjqyVPbZkUGLHZ+WVgN+gx6AxsKpoyNhojspcEAYVIkfh
myy/0rZXDRgx81vBo8j4IJjZecP/iHl/G0wN90lM60LNaQXMbUkFpm/XX4SCAezCIEHuCuQlS+vT
oPzkVmPqb8qEBr5JbEiUYuYhr8CJM/3VULG5kdEsqFlD7xz9eFFt9Qahb3ad83fsrDzsBfmpH5XX
BBSkcVmK29bmVKWlQhCIBxKfEa6k2G9Qx/UlV94ivr7VZRVhYngtdcDDCl/gBBqDiEOBg1X3IHxn
d23UlDEKrpdKSxy4bJ7Sm9txWgjdRzTimVckhDBrjjTBkzT9/uTH456cQ8rOk3fod/i1d6JYWTKE
L1Wkw6vYKAM+4qzl8z4rlizrmP7hDOhB7qhsyhafhtKls3097DaKqKT3h/LGk6zTHTxDFKOfIeM7
fSJxjI/f0iHpDh6dd6m5yzRsHJ1KmGvjrynNQu7CJIPPLcF5S9yMFK5JY5X3ZzpsuYRwCCr1vj7W
mP3VKrUtGz34+Mxtz8UE+f/HfzA9uC3uKdTQFFS0vQywtvBMwHToQOycuJoOmeIjhVJWzyAS7gxf
WNxEAzPHZNIkdCVSlG/5OiaTQzYThoifMU7UpQ0k0CADQ0t5kU3mD5j3KhuqyK3GvZyeGOAWL8gt
FnnpUAR2wPyb5Ae0X63j5mXiyIxL1Sx9oPzEp7IohPdC6OxhgCrP/M6r9028m6ligeekJbD1bgJl
wgHLreCwCpT6saxVT9JHdL6yLR23wNHH/aFCEYKwPwe6p1nPmPsWXhKJI0U5J4ibeJSNqGsOkZU3
xKsbFoQ2TrcQaZ8He7YqULZ/JltkYbhCeHWpz0xlUkdNNke5p+kDudOc1e6LD4Q8jOIZyKdInwfV
CydbazZUP2OSzC4iV0qSQNxwfCnLZWPXwTaUdpU7VAgu4vo3HN2IKOsEP1LLxCWE1FDCHNTwnjdI
7L550GRo2M+6AnDS5zdidd3juTnMd4sn1BqHbAIYSKcccPY3lHrOTPYDBccPViwAN6kOfqa0ZrDi
stfLrU6zCeTFsocozhouk5K0Uh0brmPnDcflPOQGG9PcrLui2Cg2c2lPNogIfrdV4bg1itJw/y7m
YsMqqtJPzI0jWebBwreDzA7tdHPBr8idy0Tx3ICFfVZjwM3d8HCW7Z519tBSt0ekGoLht01dek2a
q3tixKxwUNfI8/oWKSijg7UtJBWZGuAW2RBOHLwbSrfTXntaOprfe8/ESGmEbcIWxj3OqTGw3V7f
hqBXGYSxxHjsloKababBCtkPn/JaR8yQjIEVeglrHKn0V1t/kPv+CXJoSiKVv/ISoHnRIcm3IFn/
20tziEJsFZLPbIJGiP8Smlx/zFf0B0UxvxJvG2wNlssgMjLU8S1HgVJL3r27n3FNyqAYuDOdd5C+
sRJyj2ED3p9OVkbU0s6bKo0zD8Xq0aQeQt4mRJpkXkhLWx/OSAA3hSFMDCFCHTMnrM9JXQJi+D1g
fwyW0/qhzcuk5VsEC3dxwzUyBjxixt/LejNdv3Bs1qNg0FZ+py0EYQ69oQ79ughxlaSRcjHXpIhv
YAnN+ogcTd94V3tYjiqJMhpHJ3zZHNqoHCQFBlS9eDj5sx14TPcpQN4FWpu8dcpqv5/xPSGXukR0
6KklLYpZJ7T4+id+FE7xQn1TYppQD1IpqdsqAEvIyMN0Sy1WeU9Fh2/KxCKWribvTMP4Fd1RUv2X
ldxG+foG/lKhjdohtgIaGvSZ89BoESMZiFKHsarKqhKsPJlADrC0MZZyOqaps1JmpHhsZnC8tNi8
UPa2Z2yLsV+rayy3Mxvr5hqiNqEj78sTF7LgHBDks+Hshy0iOpWeN8Ef/hYws5REbTD+YEyuW8mk
EmxsrLg3Jy4+TU8miJWGmJWy8EzW1pVWn9tOX9Uglo3SZnvh/cHttS3obmO/GAlDPfbYqA0vbehy
yPF0PvztEbZG0CuoPaPtfuu2MzOIfXHZmgv2MkJbP2w4VKv8lgGMtyE/fibPJbt8VSKuK4Xp9K3n
XwH7MmK+s3ipY5yRU9CSqeUSSH1cb6AatfbvbKUIXBalFsuI41npwxW20g56tdoFHY09TKDUvoMl
snhriTvdUVAsi/YjICwKH+DQlGX1lN2zFu+OXZRMiFtKqq4isWQ3A2DSxLOYX27oaFPPyOSjVBf8
lKmrCT9lZ39CRVdyS6rYSussTwP3bvysf5tWtRMJua8whaq+UWwe+29Iek1lCd45KA06zsVEmCQx
0Ca1aNZeVaL2IRoRhXrwprFpE2Nm4NTmf0QKdveyQHLmjZNdj2XTU9uTC545W9Lq3rXhcykdK6XD
6J/BPIWUcdAEeayxtFh1oJD/7dAS14t3r3VhtpJq4/wF/IjZvPOoxd0PTScW5T9pTYXKJrYqyirk
GYz+FZhWD8u6SGFEKiNrZqChTl06HBpKUhNx5YPMLh6qsMP2fDV7i88U8wfiXS4dg2zkr0ig1YaO
TRaQtddNwYn4w7x6uFAUZIHMxLXZrLh0wysRodtdolbDY1LQR2ryDjSLtSbNt37yRvkbE0IiX2Ay
TrXAVcCDlq1rd+IDlmHynTAGWm4m2BOvjEERcZEukjmdLfWWCTWnvwiQNO86YKZNxYNvw6MjwVUa
oFGNwXoCCroqdq3VNJ2GyGOW2IRVe7ki8R08DYRN9af8LXLAHozuX9xdQlRTL0pw6toHMBPq9tIY
c62FoQMZnW2mf6cm0uxZNoBiYfXp4/lgG6tQW5rXrIcV7F1W+Kew6cpUgVlpk2mk++rsx8SYRm6j
yftB3HRQ/lmmZZRCK9mNbCbaEUL/gfhxob0LF5YCKRFtFM8bKtDuXzyv93TxVrqInXbm0eiXejpX
b96BsP4Jjeaw1kv8gUwI+Mq0RtMS5IGXpiDE9DveQGS9CdZBI/Dcyp2tKIFt+RTAK3TThbq33/J9
VEl/RHqQ37YOgqGp1odv1tEyagrNuyUqUQ99TQoorLmDOlYRP1xLsWi68Eq3K1o5lSj7b9eAbd1p
llQgI2foO0x3arJ9HkcfMHIlPKAJDhY3fsZ0WLwlcemay98KND7wG9DpFzMs0maDRBAmHEPvKNvp
PFMrAcoEXWCxqF0WuEvpsGOoHdeINbH0wLY3R8huSppUCrFajNNR9Rs26qoOumJWgFRFRhZvjyYE
hLLSLOFbBVZOEVEVxv7KjAzMGMmtkbCt49O2QYb8SE90pna5brwjeWv8dTzByHADSL4BxY6+jOEj
YNxHjjwHcZKcQmezlBe/kN1wOBjzULzzvVf6K+PWPg9xvNCPwWjSgNd7of3R3UiRzJbr9rM8dzl+
xY18VcGottEytq7IctidsKdVAlfr/eCyTCkIkEPoZLcPpZAwDoNjWp6UXKT7V9mu7emNL1+xXeEm
6QsDIwOnyhCbJ+LJN686ssZiE+GBco3rYJMDNQOwHjIKBTkmU3EJkWMuuLfp6YSGuVnmJbJJVXZU
oUwqaN3A3RzzS/FzPoLGNcUiVqDjpBcbgavRzjsF6X0ohR9Vt3AMi+B/HV0rkrYKG7O0Gl/VCYPd
znEJXNs/QhzJd1pVxjSqertxPbqWHPqBDvBphRJfNBT58Kks6zz29T969rZriX0L3DN9scC4y/Pj
wYQiDhKMgu6VChXuARpfxgfgx6cJGGvuB5OBIMRgpsoR3beogTrpSQG0OyPqMiZQNO4QzI4UQjUD
aqdIGhqxyUQwKnprTLqcGHEommFmeP1rkcoQHMmrTU5lL9ZBe4aUtmevjlYJX3qjWRobbBK92NMK
Xla4F18ga8+GZU4p2k/rygd9FA3JFHX0MB/ZE8/VBnscefGIB364Zac46tZ5OTmf37fnMuq+ebiu
634MPwY3GuuZTzsn/vLZyhCnVusLqnMitVWCHhOVmlCg6ho+NONFwSgYnt9BfVjOWiljj8CIGVya
J7zLpi83LnVTada6NYwMMCkckcYaUCXwwN3hS2mOfLc/IvGicFr8Kj4DRy8MdW5B98NaBVxFUFMY
7zLozHvlWaJvcXdOvAjCwmsOm+i3DlUFbyAe1gNgDHIVw5deRVB73fdT2TgK325hArkRzuMaWFy4
7ZojFPd9cVFMRGe3YfY1K6dxQICFrRu3PO7vOtYscn/ODYv/Q8UwIUaa/DcwEJB1xv2Gxyw0vrqu
px+ClfuiAQ0D5kKBpW/ipdupw5CMwFNiFN/eabYZFd2+yb4er9w1ydHxwcfNu6kqIHgd0BP21/WY
pR/OUsUSKQYyCzLRJTw3R1QgkOcMkkhryZC3oo6e61IZN2Je6bKYYAT3CHVA625SGi1NUbs7Sm75
edcxh7w6+o5AI3AUruM0Z/yyk0upRdyyPv59ySeoZKVXgHJUqfZHu10a21+4aje68sUyVO1K3/1G
dZGliABTw1EEXu1gqZCfE5S4HwCYn+LkMYUJVO7v8KL/quQHnuezQoM8ZzI9Uaz8WxzoG6eOU+fz
ifDe7u0EQcArVUdwVue/4S5423jkWGNJAywEg6Ir1h/a6R6hZF5ESUApWg5J0E13Z0/imtLgemMo
eWoc6JdY/zYKsRAqv2katA4xo5PBSTUruFB2smJONvOE9CSwsAUCR8dTio6f+5fpLNeRwzyoSTfW
P2NOugRxofVit0tFRw9RJc0kNtUccmiwqIEQJTB8pzIZbdUTW1M4FgLv1klz/XO4W+ThgPv8nmpI
QiVt75z5z8JrDUOKCwJaYQ5GjWGX37+cfCaVP5a5I/kZLyBfPKNFb7PYUj4N9l2ofeXrJYLOUP2h
6gc0KckJBC8VwyIi1seHg5BopvU1nDREj1Fpi+rT1a3fTIj5YhYeMmfs9adV39REn5NrWG7UUk8v
jzn7EcvImnaIHFco6rI+g7ORdY1bRCc2KXC99i9CFJ0Il6E7B3WvUKtDqQF2e9SxK/7zode4zoDc
dBom2XxMc/T6JhpH6sN0fPwOHFN7eRmT5JfVVNdMZ94yMOIdRFXdVrRy1n7SCOD3q55hpVPFhRmQ
79rbJ4XMNH6Z9caf1XJ9MTTU5kP4P8svH4QmAgvCG4lCg3ndIJ4vY9MZUwSYbFXzgGzIzC2iAyN3
V1ttWOGLXwSrJM4YXiVKhlzNdMenPF0duyl+tSikZZyZz1Ji8QLoUnMfw8WJzjXBRjzWFmUp9nvX
lHlognVYKmxGG8BF6qywtK364nR6x5SAhHtJs/gAEAn6MhrcrgObMCOq6wSRYAPuiFXIEzMzDCQV
OmGbOV4JmkHQr2b9oQJJG79QQjRceiam54pib1p1yGZ4VBSq98ygNmcuZlHSd0wm4+/HRKeNhVHu
cGIIC4130HfDG0Wv8DbRYLGNDr3AApUiovu7JwHlRyAdYuawdILJFLUK6ZiAOR7qKQgdS/sCYy3H
7+t7nP7pfwgSODMk25PP5bUlVS7Kd9hQ39P3+yOX3n2sR+//VqZTbmTV49F1tSxuf4PDSHQr97PN
5iZJnxUuB+PHUB/XtVHFu+uxhBwj5PSLly8yCcKfGfIEwgo5A1ntSDFFpVDEjO1OZj90+/ffSS20
fNd+f2y+LK9j37rC4qMvihJo4MmPc8zubK6povemlUwkmzMRBXLuavOCsqu6YRQutBXH26PNeryS
se51lP5fQFw/Q7r+RsT6uVLOWivhR73jnnk3/y6r7G9nI3NhyG/WaCmX1JfVCqQUtU/stKl4twxc
ZuIhZ7O+zBXCBngOkpZCgyXVmSVSv3aAbGXWtMWJzKant2s+Ja2fCcM/1h2pajELBV31fFXX4N2X
ehfzxfN7YjY019mv2MiLNJojjIdTPpxQEvpF+OrwqHgMpT5ULX5iOG7eqjOg7Q2HUUDCAFHGcArE
3Wj76p2M7LsZbYYFMpuX4tGHp08I60t1cRQ8U+b6apS3d2HdppoX5KwP5aS7DXkHpAH4NLprkSAA
GVwMsFaAh6RBZ+8A7KoJdzqzY4VLm0j3lbyLRwmqtPUs8J+Rd66Mspk4vpRwiVHV3zkJiy41D40L
m3H7mU3efKFld2MO2L8iz39jAoI9tJk17/h6iiO2Ff09wMJliQu8SrEeVx9w+QkwSGpD9+PtUMbA
/wxrRvwlkcLed/ISxH4iWrW7RSefMB5/R6p1r6/+j9v1czkXNBfgUveNCtlk8F+PbAdrhlBRa+JY
SzjbO0zpq2GkpXrQ3panVG4hhX7cQUmgDHWQ4kucPrR2EeC12WGqeXaA2pCUsW2vjht+GpdSNNhe
1i2w9SwExHysKYsaNYb4mQUyuZzoIMIcI4HpsJX2QxGYYRWhl4ETRb4KFpNLR02u3aUPq+fBJSoO
qJYH+Gbfs1U1FPQsnS8L4w7GC1dNwFtqK/wHsvimOG1bbJi54iy4uHAN9ZODJtGAb1asqFXlA4Zb
g4/kCcrhOB0zWXv7IJ4YnrTe7GzlYJdpZ2Ip0bEmh87gRgWHWbrnDPzz4NeDaHVlxOAyoCz6oxGk
y9uPqtHZu/RVaQrJ5Pe+fTVQ3a55QuZQASHSViPZvlFW5bGkiTuWSBunUKMLwRS1ha8iH4bevtt5
stnDrpuY4g2bwKKBKI7yLH0y7ZQJrJz4m1pNQU7v3zYfRUHVIQhRjtpobNzJmjLVCUzW/3YKyueL
5tePL+x0GmSllGdEi1zTy+ow0SicqP2GwWZ80XumidrI62TiLYW8Pm/RTcoUWT+QXGMAF9k8bCYP
PyZkj35vGzzups+Cmwij+CDmfW8r7o8y0YaGqUfRJu+ofU4vj0LDfVKz7zsIc48AnL8J/KaqKi2I
Jcl9NhFVbjjvt35m8nepVhd6fFePnMdAuxptTVqV7Cn5cT3EZ00wuZ9ncqOVkiS+ypqkOL2WBtWl
2k6U4VXGKOLyj08GZ0wemRpu4zizX2bO0x0s9ASjUM1AnsoAYpFtYf7zRDMh6TPGIXDxFOcFT01s
CVGdNUHSp3pSXGdCNivZj7WyUzXwjDC5V97z9YDkEB2aK2s9/cDa2KGlWjtdsgC2NvXkdR3DqTU9
64yWbbbhog14JSfifImfiGDclM5DLFlI2lQhaYvLDbD9DYbFbsCxI+ZB/in8qN5c242mbqChFQiT
+WqcHgf3KMZmHkciikqQ56k+FAGIuqm7/gjqbQ4+MFplDnA1bJSsP9PvnSb32VaicKz+JqBCJyqn
e0Awv3amuo2uHsyZClv0WcXrYEIg2mLSBvAKhbPaSP0MoRpGeHdJtLMmEXz0ip3HbxEMJOcGuXn8
V2iFtwikzNxDhnAiEtja+BeftIME7tm8ZEmdZ6EhSU7/qe9m5RidCAHIYvl8vYj9kUENpkdCe0DG
pfK0XCAIvAlDrDDJ5kypKi6hIccz4LG9AYpEKtd+7eVRf7rbwoA0KTRcHPqA5q0YeVCPzROwspws
6cPEuUhNxx+QSIKLCq43BJdZmU7J50gTo2LA0OJXr9UVrh34QVdr1BO+vsNiTtl/kvbSRc6vJ0mG
Qwj1hbIDQNvMJZbKg6Iu2KJWDlJRPMF3RveJ97ia1LgYlY+w8FN98Z8MG1/Cxbq2EvWj6sobBkLV
drC12KS7YO82
`protect end_protected
