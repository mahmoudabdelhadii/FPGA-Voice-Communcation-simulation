-- (C) 2001-2016 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
zMP9inTWtieuay3/j75LOJi6BSd6NDDL6J28CDpGrGUFBTmdJjBAUnyEr8t+JwDt0oV8EjLFJnB0
jFcy6SJq/nuh8ly83/d02cqFQa5Nk/03RDAT/blJad99XMC8WAgn0MW9pZwnXOesFDWZtEgitnyj
e4DFMdxxUvJlKNDnlcoaE4I2wM9gCuXIz153R9Zwfws3HnpJTZlURxTIfi4WF0bg13fJ5H4+SdJr
DC44htnCZBpDsKtlTK8Ujv8cKwOz/2ZvdVQQ8enpMIPpDBLdnuz4mJE09LjfuPAT8L9Roleo1cCk
smVv7tp1jUuBzZTGKV3a/qV6EJFdymdNAdx2iA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 13744)
`protect data_block
IXy41rNPBBxe+WWBLT80JdgnSgqguZlAMIFftgtqNiO+DyHTzlwltWa0jNYMMcDxoGc0qMDb075g
5acuwbzJttpKXXZsTQy6jUaNXSFJrWDL+kd2zHTgp67SayiSG50hNzGGBc2guGVQuF7RJzHcGdb2
JR2x3gRgfWFKvn72StV2u7KhcsYim5RG8dvN0h7q/hob6M2ZytQ0j9Q5BquwZR+ZZBCxuw6kuQl7
Nl9hzkBZ6tdnqdLGK4pJzFXtgVKoZMzFE7bkkPR8MQAmEzZOmSFUJFKnu/Aqlo4r/N5LIGZVA3aE
hBjz6hyCdEB/sLb/juBKxYdvrpJuTzKmWETkcC9dg4MMOgsl2L7Bh/LUYCqtQrEBA+Jrkht3izop
oAEVpI0DtsIdt1IfQoYI1cr49MIGMmSUU0EsewCi+UTYKQfvUdG3W+dqgnDPrqNXwTrjaNfRC6z6
XJsicDeKEUiNGcCWtr8OSvA6jsuAT/oj8BDKTMN43aWhuW2lw4NuscLi35jsT7TVTJDML/n76Yk3
J2oXTMnfRGVFI3V3YnEzehYKZepCgpBDY+0BxMjVj6eSnPgbDaTGDvm0G7SohWv2CH4RZ4Rv79RK
aIRn47gawUcTbZUpp5mkKUpz/nB38/AxPurEWeACXg8+ebh4M4mKIVRpNRwy2PZ8GUUixG5reD+U
7Ns41IITym9BpmoKK0lNBYPfwSRbGRZlsokvWXEr343m3ng/zLeV8PTtJXk2cDX8Ka99gW/AGKBK
YC4WXQ4aGInsyR3+XNgbTjLHyUY/qeO3J1ZkXB3FkZ0v5A2qRHuCXwcrlW0LJePLOFjORaxTxkaj
cwxQ+Sym1Rvyf5oaZotLboM8e/T2ghvq/iHtDBeb4EctVibSedBvQHIOb9wqYxJoU98PvqyVIPIy
RozfxJneZWH1ySJrOKbh5Bmehg/ZmDlbFS9M7mqphHRCy0mE8NGA9GzuFGZ66wCuGbjwq47iTrZv
Uey4tXJHDh9bCPcT9GcuAyS4uA7Nvb6NgQpjk9YfQXNX1F0jXT1eYnOcQHOEMj0tY2fLz06jSj30
upGzOhi520KE3MJshYEU5FJQBSyAcNf/SvbzKv/HoB2ham9EMo0oJc7t1FpP/ShkwvvrmtLtbBGe
sh395MOlGFVs4Q7cK1bE+D5oq9d0KXwsTfxk5r/QIfppP4BB9hUEESm2/QGR2Qzm0hNYVZImko0R
crhY/j7m5pulYwQXse74I06wCKe2bFsxZaQWGhZmd4sMp1fz7QDh+lEcQSr2xEKX8bo7o4kob4Bb
Q0sxaQKfIkg1a/gplxkCCr2LEyJB7oE/EoEjzcaCBfrNG9o7xCx3iRBwFI/SoTlSBN/DyDJlhEhi
r0vMoP6rQtrV2dO/K5MAdULrCK4HPk8VhNSh6ZME5xcPVeFHmItVuSW4hET+E+RiZGrkmFL37Ahc
jZuE1fxwv/i7ooSHzO7q/qEr8U8Eg2x4moidU4g7Ke/XtmQp/vc8p2lscf9MV6ZYHXo/sAyccl3X
I4ggO4BXNT5B4Wh8TgIYmMCMGTWgy46X2PoVDAuaYeubDEeCWYjj5gQbjcUWGak5GHbg8W26lX/g
H66xQCuBw9OjRj1ceBLOGskd8aVKj6z5dG1u+P96sjVvKChroE2Bx0AJrvaYednmio3X7qrJmfqr
rENifzSHzHPCSg6g0ZkJo4iM+5xr4frXXZ5F/WR59ZIYgeOn5PqPsETb6GUZsSKBtzARqqqKvzuY
4XX+/cEf+yelwEfBUNbJsmG6OkL5YhDZMjtuy7oLZ07y9/kl6UTgZHUp5VGDsqVtZIvneisJ7jJp
Y1Zb69s4z4BeBhb22m0oAmvjTx2pbDqWLGWozyq72ZnUzFqWgy4k0LgA/6zM4e1v4yKU2iB44i4Z
eS3QCikOps+V3n/aDfYQONNpwgWSMNe8JeqCIGnXFAtEhRxVvMVKzRE/LKtG+se5t7tuqOjZVuOU
TT/y/qjJQXQnJ2FXxS6niZcQqJDs+WiXmTSzF6ouc53J9YsBmC3Zhp1wHn59yc41lY78ybyAGNfN
rC4csnJznzcGWdUAjaMJDnPh/k+Xl1zniSN5KsIdn+8yPJCc0GSsHagI4GvWNyGqrXI351ju4zec
OJ0GrYieXF5hDQhBHxfZ3WsQdCJHEYaa5LDnl1fN+fpwWH56qObhI0TMO99OGhSaPHGNrXQ8QCvP
BI2BEB8LhP0/Gji9KtPbl9VIIJG/xelrz5GchJZEksU44IFVPfcDm4n2dciEZPBf+QBCI00lsQ18
gU0c7D+stSHyHB0QqNn/W1d+p9L5xssEtxPGkL9GkJWmepNl6mUpE77NxAU8RHnnpgr7IwqIQetA
wDyOu6lJv/szJFj9AqP3Oc/z6NFJysz5MN5hFgOWcIBkfkF740NOysg56LDynjaWAiO68yRXBZ0A
IFXOURVDKuGUNUQkkWef2xXBbdD0ud/ERv/uduTc2DrM1vhFpNbAdpoKyNvF6gpuNwFwldJlt0os
m3Aj8U7fCCpOai2MZ6j/bUs7Upn9nqesebT3RNf8KUZCQ1pq/jsEsCRqgXUZSAfo3m/vo+KOw96I
Ep+IAw1wEG8qg7onlK94u53YbBlpWNiJyD5LYcHRXOeXKIS8HqfOhXl1h0yvoInof+QlEHWdn30L
SPeYWFldtzXQvNC0C0sQvtnImruTgCDGI84kHwd1UjrvZXufhqd/mSek5GgQ2ZsQw/yHfjebN7nQ
YsxwFRzws9Nmr69pjVk+FpUyxVhaKBjJLFORpWqIL32nCbGm39XvgKSPJtNFmAa8x7uhGqrMq81F
JrLxE1Zb7QaRjGR3sq473+GBxF4Xg6c5bWDN3zTZoq1S9BneEarlMTc12n4OgdhggT0Rxbq6kdjD
Btfn1Ha2ZJdxKGQ3zDablNULmgZP1hofs/qtS3RrTJ/sgEQoBWlr3i8b+RwkcXApZ40f+5/Nr39h
q3Xq6yl+u928AXY2m8s2s8czM7qmsETtpo9KScS7gR1ptkEvej4ag3jQS97XW2ItaOdu/81MLJ0U
uG7vD2bmqKHgr672f7ffD0UqIp1w95CivyaZoyIiSXWnKVZi80mNhsJBUKJcbyoK4QLvJU1IyRdq
emVhLgzSUmifNBDqLSOoKMP9ou+MPoFDJ2+5SGT3z1G9wGM08ih5IPVQ6s6t6LjzAPbHhuXH2lLN
HOmdjql1Gcg1oSANwp5861GM4MW1MXLi0LXLyd5sa4repEqQvJbKFkagK6eL0w9WX1nrfdEtTUTQ
1+JNIkLZt02W/685jA/JG0zX94Sw74aaGbbv9goXwJqQ12OOAV6ND0MVRNMGM+LgQ6i+g9F8Z2cg
qegEZJchXlShltrzflFLOwf6dTbplKDRr4VLOOYOxjcV3tYKCaEztGlZEpW7tNto8eh0LqLiUR8l
UaBXPzpnKsLmNvXKSobTZSsIz30Rz0JRTM2mXOvrHWhX8rYEGb+XHLuqZQwXTPOtA3IyrZEod+pW
M+kBkREQnK2BtLcjsK0amRehNnHZUbJJdlJkE44yRK2YsNhnicbEbFqfAxHPeFQjQB2SXsQS16BH
6mf+4ZkajQlSTiznDrFQcyRDCXfsomlBzmj9+EHKzSM4B0uBP1C3YB3aK/alxq9JDoHAEMJi6K/w
daa1ZVC8HprV1aWr73jqBUwtntmsoJaf6J2DDx2nVc4A4sI9zYJWrgkKLE+WBFPj2ZErAogJ8E19
dUmCFdiygt788D3OyHUmGsIuP7gcSiPohfGiQ6N3FxHQGcYNO1+xlkdheLKkCkuCAJJ5hI176vAe
J0noMf9SoCz73I7e+bOYFSdE6lqEw61O/ja7Pxm96C6IG5AzyyU3nTVMdlK9LoiLWHFI4Ko9We5H
AmNroBfgV2hzYyu1JtvWwsS1qPpc6gm48mm20PuFAzAu+RwGPxA+dSK/qBgRdKcT0WqbKaFiGTXr
1+fNxeKUhd1Rzp3ycSFBEeqkUdx3IrouP73Se+pTDcfeF15IbOyuPXlU7qMLmp+gIJkPqzAA5UMt
eFTmIWetwwl14VQzpDdR8U4B/HhF42wi5Qo2fjP2MYKWgxSUbxh0hrfmPv8cvsoKfRwENFPYrKfE
00Nu+lUPQuLVhidLDm777lI/SGDl3l7i0QhjCm2O1NJ5KPQSFrdfrL6QBk8Uf4XOSn3fetmie5Sp
iSncvZuY32VsJ3A+i9qjcV6vRzKBDozzVXHw9K5Hwg54644AYfs+uu0a2cLuTCV+dJjTLKKK8a4Y
h1XGVWOO4pBHG+N/cHGlncX16exLkuVjV8iZNYKyMSN6HlbkW0T1hL5fuFNbsJ0fcxwdnh11BNUq
J1oc9svdVqEuiw1f75mg3LTwKiGXoWauuulyDovA54BuDZyMs+BP0voxHY/xF4h8lBO6VfsNuils
/7a+ov1FEOzsH0sbVR61uoA65uL0ZPVa1MypxuGqjsF9U7ljYUvfBE54cfgICxkP5lMTEkZe1I+U
4ifOQ0tcZSbiEygQ5ksmYGbpkCwX6a9M8Q0adLopaRj7bn+iYI5MCfXxePZQGgED0U2f74vGxrXw
R3isdIQ4b4fKBSSPp+R9zbwQ5v6wmApM2+06fA5OIuI995ORhCwyB9XqfYj5CjA4bMj54Ljvtyxw
01BZ6lAdu5Esixj1WaFrLU1ljlqcgNyn/0rC39QPOWSLauDl4fxCjCUwplBh2zXMMMcqvOVgIgfv
eCEBuLAEGqgiVLaMU6ZEC/SzIXV9jQe2K7rqE2PF5dIOAr2GDHEUC+YfOD8XOBaXmCYU81w+dTJx
o1u4LUZROCqH1wz1naFbirp7RM48JitD9WlYlsyFt0ZN6ZaqYC/UoTrTGPHr+J8dy+Gk+fpB259K
XNwQo6mHLM4nlO5XVB9i3cAPxxWENjZn/8/n/kFqoL5QUrMTAJ3q+8D/Mqfa6+Y0CRXdD4+l2RS0
m6U5HKMtlpxzFbXht/baKFWZb5Q1T+8TQ8ya9zJIdRPE966yned+S6EytoDKDVYGIxtBXLtY6dB8
nOa6o+QiiZOEBT6/Or6kJTGVQDpOj3bN/H1gJdeAVDDOVWkQhdmdLREH6QeKbqc41yFbGo1CwPqz
5eKSZLhxclJp2tJguYj83/0/WfKJTusTGVtKiIB2WePrnDN8tRaH07jHtjDpte8h5k0guXgRp1k1
TpgxrhtHKwS4lNvDwFTF1o9ygBmipEYIol0A0qxIXpRp66JCcrha93g6MKadsSKtUjWlijbtCHyg
2nwBvf2riwkkCrNFbsDQad5GCpcMJdFHxYuTDoZFkzFfLAxPoRV9uRGaMrGQTjMh0glwH/lQfd3F
gDOCs7zoUQ+qcxiZ3uF1G+VJXS5uUqDanZ5rDq1SlGLmb0hqoz+3C+nrz7jyvJmCYot1UbOCn+5t
RdCO2+wHz46Mk/sbKwzUJQhJ7ovf5phTBjTUa2zst20lHAt4sKnuwhsWYQsoWnsHDTSMLczgkBp/
bAz46k5CdhQ/umfIhG/hspJ//hJUxXPN3/AhbE/HfoP2o+sZeNIR4CVKfvGL7CeSDR3xrfovR8Ui
Es4uQEJkSGzks2hYQ9VHYKttma31YcWG+TpD2IVz0ycjBeJg9rAE8+k0NQkQQIZXlsQHRJBSVqzZ
cYqTADdgqdeoJVzTWKKwE7Y+r63zrQLDoc3M4Vr09vnHJEqFQ3DWY+UC/j3BkY1gO1rXR4wXGxxd
OP27GWE7av8hQJJZjK+24AhV3/eJ07zZlSEd1baILs31Ar5xBB9T3EBWmqklh8d3B9kEex76ysFi
NiZLbZ6gDelHa0M1/eByrOraV6v93lb3+GXh/TrYOhWFH9oFkzHH0ihdnoHMxND7es/7HWBWkLKq
U5MEuUzrIvEtt5WaslEB2exAjEeB29NGCWUoIBGwgPBegChCY27Ti61tA8rvfBjbBq/BiK1HiHr1
yAvMIQ5tnIeK9lwhBR7BHooE0g6jTaPylR8sQOh1tdI6aWDgUm/j2Qz6ECojl6kPCMauCflZEGR+
v+DlX9+AvW6YF4p8pk+hJL4Tva02p/5VEzTTS4/AK8sgEFAc9xMa3ljfuKFacV27aPnxU/PySuna
pbv8h0NiPm6iV14WwD4bg9JNG1wyhwM+dNATS/8kNn+crcsKnUlC3nNO5y4phx350EAihdFlLdHA
ViNQptHoVWOF9pBTotQeZoa5pYNk1e1c3BejIT2s5wCHvnH7DjcSTDaVphZMEjPW/wWQUFZRsB8i
Ig1kUqE/vpLpIZjiPyqvMXS+hKPPkrn03T4Ctzephvs3OaljTIjjYZ6vIEL+hhbehwTbPY+z8yBR
Y5gzfRlk1jBO4YOObiPybNwbZnZDd+feVhlxIJ0TQl9JKID6bA3TaPxlGhGj+4ofJimzXT+c7ZPy
RNexQbLJOJQ5Hhix12Q31WHtz8d8M27FhC4hTIWhi4VKXhN5Q2pzhTegD9d+JwkJeGK/6E77Zfmz
Al64yQFx0iSjn87l6m3HysDWTAzQaiaED3EdgjBttSjtw/pVERO6GMtxx/BYFnisQn1Ak7QC+xCB
8WI/9DfrYMV7vppeyZ3tj/VpyzYGN4H2JU68YM7ySt+m7gPvo50P6rEIJk9FkbioFsv8o8Fp0nw7
sCs6ML/4Tzt8Bg585RvnMD3eb1L/fCJKeVX21cDbtli1N/3+UysVYiMQW35GLxXZOIo8Ewf0kckv
owA3PBmUQunqd8LpeoIzCMTi6d5//Til7tT8dmonSIGT9j8WqgtCd66Ds0OLRkqJ2ypCCUUfOYoE
T+h4ewEfoJp3BoVro/w7/hoqWmH11CA7ecJ1rRXxwizy8KSzFtsXmTLibK0pmmvMR+MbXKbMfXs2
NABpMPIIAQB11Xw4tMpLc9+IxamustngMWQJO8qTrqpA+ks4QBwzG1ABfp6DE4wbf3A9uAd6VlCO
Fg5VUL1sINLc0T3GTso0fp+/vBE67uA6Q0fJb3PEctFwPM4zb2FWu3lwU2EWh7ZgVrMIiNAjvJmy
16F+unoSRNKJA0ZKbVpU7BzSwzgSqcaqXAF7XroDrtqoHjatk9Rnl1pxfcagCEc/BgTZOIHf1PHJ
AKWy7io1qjLyRRGx4p3H03dXN8mY++pdozPJn7lyseMz/ZYHNloenFhpvbXpQcoGf4ilS3VFRQup
a55oz6SNtPY2MH5l6vc5dGnTQrUt1Nt46FQaOFQKoRBoONIOHTBe2SjVxFKEIksUGrS1UDapR837
2ttbhtlgXYFS/ehKt0Xswr0gv9uslREfMh9NNaAozf5bwhW54Lg4UIYinL5Cf1DnxA36HsnaXHV/
TpD4GwOYRMqdkX7hZ5eInfQ1VASeHD+wsuNdqPwg68PZp+J8a4N/GWVopQGoMfEPzXK9tAvIBHYf
s8uPkFd5oJxoa5Q2qlYOvdt8Bq3/r84i22pcMZXmWx+Ebn5EZnv4bwpnI5oaIPeih3FTlBvo9mIN
fKVK12VAXRksEZsVPWYH9tNO2WtVUNJ/UdS+L+E3243oWQDRtS1hW9kh/LxUjaZx/FoBI0NFnO1z
OInOCGwhreUtR0Ikvskq3xX0qqorHxE3SCebp99wmWNSICj+2LthO1NCvW0XsiYFLTaD7Jc6lkV9
Ru+vY+FLX1PaftNxUwGdTLhgwyVyMQMZZ1hRPZ4OFhPYJQ2BJNd+NCetqUtRt9pcBrX58W7oJb08
pg5BzuQgtmP84YN4/aveR7GCIJIGa0u/ySsUcn4+zyM0/xASV1Hpzhpraw29fKm7KtGyiPANQOAs
9iJwUdIgGDEFaudGc5C8ehpUjfwPKja4EuBv+ctRpSmJSydx5VYXmC6c6M3fJuqGgga9i6Jd+UrF
xnBZ3s/G8Eirol+l80b/fnZWQAXVxmTo0W83KTrA2RywpkkXOSQSeXVooPsm5Pa63eKMlboomeXg
r7gYBnyscrmLVoElsrulWBxg1LChpInyN4kMSNPPyEJOYj+a+VnEiL/QTj3bshQYueAlXRZci6lJ
Z4hYqLKuG7PRVdrhZzOUpD0Cp9zDmc8GerGaOzxTXOEY2PBWUSIz7alCZzuv8GK+CKJ/KuojEc+R
HmkLq3KSMrba6KgPtuKGbHKoCgXPRkpzSxDjDJ7TuUkpdsiM9FzL64jhmTYtoCSNsawP0S4lqBDZ
yABKyv76kYz9Vvc+Y5QPRISjh2qktokMGFwnE2r0IalllOQqSrOIBK/sDKbEDNyjTfQj3CX5oHXE
vTAvWDXNES9ZHacIFc1RHp0IHGsJ3HVACrU2PHcpgjVcxOfuF2z2ilpKZaLb+TWJEYJGF/H6kgDV
ubdFquFEXtSbzNp0nUShvlecH1lRSaTERuCTo7Wzvscf7mD8atkctUQ8UqyPNQDLietjDyJi2Y9V
dt09ND3DeguteMJU3XBXQb5xnehaimX2Xi434fbmMqHH9dpLEgZKtnuqwjt5e+aFZ4LMuSjKlHzz
kiBhoGaqf2r/tWrs/df8vutb+2l0PfE3XoKRi7jzBWAL4TMisM+8FI71R2OnftOYqsFuoKyGmV6C
dzNgp7lFiTTycDz6EeBgU1SR/9Y4/EOc0efx2lC3VHwhrC05W889xhuCp4QWRZa9liT69xeArUJs
WazAMHpepTBgrROJdH+9JnipEMNyk2ZI25ptrC9oIALdruXcUsKGgYK2XLFINiFGKTKetOWEnRaZ
FL5YigbOMRJDD0zP8VBL2MAkTckUDNc+HWh8s/kYgHXKkqmsYhyZzjEkXNFe/y8jw8IEgiln2Dye
pisv5/QsxkS9KmYbvZG/KsQblAeCS0ZZiVGtGqKlNPoUmDYXmTsGzaWFKjB2SwDSOg69OGRMk+El
3zGVrre6N0Aagfpq3c8tcxJumJRkfRngPiaIzDedbFQh1zrlmkh2hRnBsvwxDy5WKupSQan1V8Xm
ZeX6J6MZA3aZNBIddHwhEkSGOh5jp4FpA0HBbQnY0/KUCANCx9824L7nKZTkUBOTSpMn6ZTVlu3H
vmpsZcP3DDd8l2qQgBZd+wqE5RIptwheHSF4GLJl4tthVXny1j9xY793ai17wdtrgbWZqrGrRjq/
IqUIUFnpPqukIElKERwYYxdW5i5k/gsSpZyftv1pH9hCVFkaLrhzMFtybuI5pp5My5uDRRY5Dp+G
wmyclbLjogxr8FbjjNSD1KHOxXHJO3kOhUsY0K/iS0078shIkBXITYoJArwagJN7zBG+MOqU8DUs
7/umeEVbJc0PQEJ/iH/17CzsQWM30/t2ViqL/6Q3Gc7ZMStedIHbGBlBLet352HkmZ3v576iz/ic
kHlAG5g3ykOGMr4Y1FhNADovWeYCua4cptAZzg2YGWN4vux2o9qBaKAda6cTiy6Sb9z5P75kzS2b
H9yj/UNSJo4OjodX8AXSmB2owYkw5XAau+7JrozUWD6+TFKWdmSrGq0TDQwUcdfhgEBrNEEFkHhS
Ea5IiSIXvW95m5mesTUwJo/ukT9evHVSphd1VSAJtgMpoeZ2CYKzN9lUWiKbpXISjz27oZJWteyZ
3Wx7sgV0DJKmBL1bOks4u1MeRL8D9SK3WEbocXYJEGWdej4KH2t1bsdZb4uslTpkNS6uYvN/BOGK
UvkLy+lHyKmbzZoRPifj5bEuA39gv/NtBd3wDeCOWxMshrIfWcBMjwyU/ciC8iBJ2jvaMVxz74yS
MqiEA6DgNqRXBtNsngLLrpyIXM0B6kWwlPMV02SO0B7H+RE0kwHhcxyvtho4asTDIemlftVVU/Qf
kBknSL2n03KLk6etJVP9+ofep+bmpDMnkc6EsPbdZN75LVDpF8aBDRt/Ou/ZMXfso/2glVcwUCcO
p1ipc2LhtEDZDcBWm6whuFed3r6T2TZjRL2MLp8JJAVzXowideBsFUPuIxOs+2USomuqMKZbklqu
oGDvpqPVvE032tpt8Gs9pJq3Je9ZBGVHMN41Zhn+0qpQk3nJRbSEkYV7EQ1IQVcHJ99RMIxE/EWH
2phlIDL73eecv5ndqm+Y7AFC99btjwlnj3i0lhC5SFmJvlP47IGaU1NESPNj2OR9E9jF520TYk5K
eeg+32fBjqtaX8aClAbF4a2Fm5VvqxKMS3d6wqDKDhaclRGkb8Z0KGuiEsV5Z9y7iz3Vq5/gDHp6
W8VJwhi7HasF0KJh2Am1rN5rUmnSWuw0pO0o6grh7/bdReyH84NIRYMnIEmtg/BMoJHlUGpWkqlk
3wpqHb6OjwMnV9dJXEdAT6s/itxgsJNf4zddre5KZMIQrcSKQj1vkbKapx/Cy9+q/K+6IvQZOOjz
NnuHKqAGdxurODgsW61VaKTbO9STbRKIRdeCHb/uJH2HYouRlRfqeSqBnPHnIvngNGtE+V0lTDyE
aKuV3NF+fSSXjPZHArx2gRRCuIdOua6xFZuOrLWwdkGA0026BPcfGXy2q2qORfFOWoPq8VkBZqml
2+JHFyp9cr8jARKUOlfEmom3L+A7opN+JWMKdCTa++VzMlW2UBiaKWSDuiI3OfP3CSlij9R+DHUu
ru5QEvMuBnX7kj/tGrwaPQ2HOUix/uPUHCV0LHg2fdtIxiRn/yaeHkSFOSGDgC2Z7KbHgBV+MWCd
rp0/aGmaRf+g86TGwK/H6h3gQE355RY3Fx9edTGFsIlumquQJDibQAYI5N5QoIJSjp+NOWe/Jnj5
b2fMuyeD3W90pOFBtNHq8h8hZdrdz842Dg/B3C5/ZizFGbLYiPMbC5jAHqivH9IlsYXGKvxP0U3e
aaWbgg4GJoF6NpAIcNz1J+xs/gRLEqbk6W1AOcUW1QaovoXfBZQxp+o0NdIiXWKyFzHU6p4h3ZAV
luyt9jxvncVHsAaCfdDqUqBTF/TxiYY2yaSi1L6ZY4qjB62E+xD78YuGscOrn8+o9x+y5psvXppG
IUioNf4ygLD7sqsZy9nqzqtP/evDcz5kBAZBLUTU6AyCn4MrI9smmhYoKXAVTi7QGqDfcHfymn2A
oA+nseDV6ZVrX+JSb1NITr3LuUY9kPhKPuQiBFXmqAOucUgVP6ZIVqf5jt1sTkkzyJSjKmxaAU/+
YvAG9WJJqxr54jc4EkqIQiV7zBJ4qwlOY6PST1k1ir9nG/YOb+SmtQlQhB98D/obPaVvQURFOW5m
T8Pgeb0HAuhEvXsgTFiU/J+IPxB1kJzKBOa2X8k2Ap4evrBz3Mul4b0cJJxkBQcJeTwSUMldF2rM
Ne5LJpmjzDbl5XF+o+YtV3kQEeoa0m1ptbNbxKMcDP+0Cs0etl26cSWp1IW5b9AzokilXJG7qBOk
pjnvNaZ/ER6jO5tfQlQxPMQD5x287ZgalPn2odk/d43EAfvSqW+Alin8aXCm7a5+LWPG+jSH2ixn
/JZl4DOn2Gy78UKAqNPunjDlfWTYpVUImRaIqOthceSnW9jKYqtZd3yEFMD7qAtFUtLvCzdf9UXf
sf4YfS35EMlpdR5XhLG1epWq4B/scMRKOTlZHQ3dSSdM/VCwlU2Wxm7dBnDF+7H0QLNECznEo0XS
pkbx3sQsbi4TBDESgxh3WwvrsId9U/nec4DA+GK+d2ejSKLnt8RnAmJPY7GGfOKwFyybg5Phz4hf
nDlVPWkpGAQmP114B8UQ7b6GipqqqXIA/ZJiQ3CuAbnCWKFJrD/BTZONIoT6zWRYfAwO60k/o51U
hJ/wsehb+DT8B4/Ye1cDOMfLuWmq/ypZjfmKU/STprR868S5+QRgdFCd1qfNHZpUSRQnDC7e2hlA
ejBHyl52fHHVPEvqLJiPkk7JphrT4kC1d/ljozI8IikqDVt/qti4F+sgARNuuS6gZE7WNluj/8IV
KgzdIZG6KNBe+JUtJDKYRXidf8rJR2hcl+34Rb6yOOuPjHZiTJr+4CDV/Wax9ngeNcn3/f0yDNRp
tau0BMYXQTT7uHMMQQxt3zj65tViyl3m4gIl1Qt5mYaFdCaO5IWsFBEaVBC88871TKWste8LeCA6
mJpmgrTjuUuP4DsPGsQBTDKuct3303sygF4DJfzLNLJVhBgfz5IUawUvtdlNHjACY90vYKPd0pDq
W8iFcGWx8gRBzPgREl+rbPvoEqrBSELYwDz2BkV0CwqBXknXESAW1kywomIpCW37dLkfdjAaHKhp
XwgktoE48Cj4m3QDa1Mq+nk/yuGRaBTPvrmS57BjS4pRLKx21Ha6pUccDZryO+jq8+7rBTbJTdOk
K8qPdzX9YNlWtbybFijl0oRvtekUCiXaSSR5NvGCKl5oPEoznxGqq+hMoEnVQYzby75b7Mh/UAqQ
SaZFg+nvd/h2VPIDHZCPGvyAnDvbpjQUUJ5AY3Crg8yqmB7x1SNPp5oUQBapnJbjegA+5cTlwqlo
zDIhZw7LDmCbKUt9h3Y54nM6MFMOG1ZX6uHDMJovuG+NTj2bgDGKBg2hPtVNzgjeH0iIYl3pBGm9
IBmm+aVc3N4C/w5QFdD/B4ZvPTlR7mz10DX51rJv3mZqvO7xQBQn2vOqj7PP8xynYR2X3pMrcLWa
O+VSPc+TM63s8qOUyOYaQ2XixxqEINeWcbI0+exDMtVdXug7tXQ4KpltJTuEMZeO34i05B5gWIPF
UDV1dfkNf5onoVsGovtmiwQyb3MSb0+mqNTn8m3AaUqmycbEzvjYHf1RiiQUtPl54+TL/Zj5eLW2
9tfD/fWvWOCAZzjtiG2LYa0hWGEkvmKHdyRgtO13Cioi7lhOqsCGYXhP49qGaRVkPHM/WKNx+i11
brfTt82wtH29Kww7UllLOaKwhAOq5Gy4gRg+3bHY5KLqxJHf5LFRK1gu7dV4Z5/CsYqFwIE8atSZ
kC0BdKpwwGxBO10f18+utad4xswK7CDfj31SmHwqZecSYz7bYQ7GL9+V6JEI/Q/K878+GefVTD02
gtjB8GqlVE83HkgRcCtTwhzIxSC16JZtJ/WPFfg2TzSrejBcHwCPqkVl5gAJQb68CAIz5q3EnbpG
fglaW3WeTHKJ+hg7QQiZLvHxNcf2/4DMPpZ88N2vNfonGKiWNhQ6DHSWhcBe6Xhpy/IK+xTxkNhc
5BsQPFAKKoaHXr+cZEH6Eo7STrwqOsDpGxjbnje0/v4OO6vvoNyWPRXdzdG0hDMHfUd3YTL9wlr2
XT5GmLYGzt5rCsAAm8fu28h8XiRDrN+p2CPsVyLYHqG2IuC/QN9PI9me9T275wrZBk8qEjVK8VGw
Sr8qFk9RBnNDQ7SsCgdNUSCcxu6wi9uDgg/clIVSUmyRvB9R58bgouuv/4TRk+AxHCKwFhmWB2JG
3xttCiA1fL5ulvHdrRJW+9RxHetHefWd4nbZOucmWkWIVYdusNYL1jS1fmPbJ4vLn4wea6Uek2cD
SN6NtD3iVFmx8g8hIpbWjlc/u55iDVNNzhNXSoLLoz1J6Lt5A1nOHmlCtt26E5zbuLHKuxbUoQm5
1FH9IgCs85ckKopCjLZxw1AzxJZYGFAx7lSQg32vly4o3BonrcJ9ta9TTsnZ2i9jr+qSHxqsMmDN
QQGPDcKKNlnuIda9IpYQiMEA8hR/vfv3LmTsr9Bp1AgEtoTEQPpYnuTD+rtPD9aKLl9f+5pQFG7L
JG2rquvVQ5f5CP+PWCcvQMDg+6R99yHhVhaczvxqRtpdJ4BfT4MpGEoct4cIcoau6DPc/UcZybxv
+jcNMv5XDcmdd4E4/BUTiPjBFCBQ6fSG9DXkRmcTJXVENJPskGBTJ4/0Vs83u0asNKnTfv+58/rI
BwBt575rUXHAf+7ENmypF13zV/L+ijnwfSHXd0s4Iv2336G4E2KzhQ2B2Zs7k/S89956TFQK5bLq
7PEgbu50PKn3NPXGecwZy1t6lkly0hGTq7WVa3ZjTorS70SOQGe+VoiXnOeJbQkljr0FIvZ/Phzo
GneClX1qYuJ2tAxmw2op6ds06rGtfy2isN9202wMsVphpzcHRWZvx/DdMQHHErvdr5WwsyNwYm4q
YDoINFrKL2BXZkVWSTiNKH+ze4Yp6kwfAQtcyEikqfEH9Q0Oy/3256XcKv9A0kkxg+J3Gvo1Phve
KF1rH1syMbA7RP50+iyyRRVHkSt0KJEML9jalDYk1xTePd9LpUIxHHQ2Yx3lwhttL/ZYwcgX5Qzz
PC7BZukuIup3ZHjI5U2lrL63ol/8ZQp5x45N9fQBxPm89aQ7ZMl+YLQGehP5rnGjMjqrfqzr/PhT
zCy9E8JvXTHgcNlYcd+rDmV0fZHh69UkAafrnob1JothgLnxFaxgzwyhdlfx6VIk/DG5Imu8r+NK
T6GMf9Q511u9IolY5MIwhc7kBJKJibwK7Nm8mVbL0DO7CJdH27OmKSvgBE0mfiplsRKuRoT1LYsF
3w0G5+TFa2hsA0Njjumu2u2wK09jnU6T9EV2HdFQCU+1/ZiqzzClyEcbpxa0uWGw1tFkUh7zXOuu
5rOOFfkDkMDrIWVxzTeHerAuLraVRbU56ax3WCzqXZd1NrBLhq/MgTLbYXvigjxM3jlmO/5IFZqI
j0DkfoIiK3ny3HrCY2DiThbHW4C4nDWrEvDpLxD6MpMM2nF4pbSOWDvPNcbd2R7sxBQFjPg110++
yuVwMgH4/lmiAv69/Zx/lezM7dMa08tb9rG3SdBGaooQiB3v90KeAC/XNbeBE2iKPXvOt0OFobt1
SbLZ1oUq1RI1zXYDqjtjCCckHThX7rDJ/qMKqcCOysvbTlQwUwQulB/W7Z6bhaP/K9gI9IzIJA12
fHuzaTlDfhjARmfH7x7boTdhQjIfrRjCBtoBp9Wx5ZuKZ9pBtmX6P022X2lu1V33HLvIyEO42A8m
KKA33D7mCFxEQ18O4JonafNoHKGOFvcLPzSOQdnVyElh7SfZOd9S7IHtyadAGS1cCoyu901uzlgc
X6XADASX2hjvv0Us1h/44G0QdmY1Gvr2oirL6nEQFAd4ZA7r1C8F9BVN8u//UbAgOr592cEy3KB4
HfVxQ+15ymMHZ4W952DCYg4H5E/xX2ykSir2BtbhtEN7OpxUgkBiNnwhjkzNHgIOlF8cUELzmX3C
kriJ0T+3LJvjCUD8MQBusq5ndM+IvmjOwaUpc4TYq64zH7z2qthms5yLVIzx6fBvg75pY4FCpxXc
7oDG1j/Gb8EcDT78c6s5HlZqmWNHBwOTk6PSjXEulhULFKY7xiT4gA3HL3HRBUYvHlnGWMo7eB2E
GSh7KfXUePoSeOo4faBmdplVJjcaMb1+AlSssQzmubs0kvu01hp1+yAJ1PfjXC3mp1KDHetlhJBT
DdyQQ52u7dYj7tNSmOH+ZN3E5J/de0+UAOUa3pH1Xw3J8NMYaeTRpV2afNYRQczZMrzST3ftA37h
DmRmIbelQdxv6Bif8dlROLeHb4ElUl3zzZfWPUIIneAoqkK8gGfGBBK2u25Qx4y3fG+UJMYHXl3Z
/CbLGaeFkPLgrd3KlpOnuYla86g8m5mG8m3jrHcGiuBEW0B7hkRRo5/bHBk2Axk6gYj2H00Ci0KP
n2A8EYTZC7CkMNHprP7ZQRNN4va7pcGS0U4LGOeWcx8z2+83FXvmT1Q8gW0iMcFsVWrBLcILwIF9
0x8XeJKLOhbZBUD1GwPI9iYFOnWe1s2dKcxOlvYFw2/ZjtWGdnqncHAo/lJVqA4N2I6R4qRoYEL6
tu5BqXk1Mprh5/aqFNYeor6REmVzbyewqtDUTmcstoJ8SstEGFfJ8livefpNszF1rWhWaNt1k+LT
HJmK38UIpYlpTEqMJvWGkzcCp0VYCcrJ42XN+HpNlLd8RH/I4UxGZV+oWHXUvb5QpIwhjcKPwWgZ
NgRC3DNaSaloKz0NbYGKIMo+Qoh3XHnzIOfmG48xRHcL5b9Ae1jNHz0ATljK0+Mw8RDLlXUJh1zU
Bma9+JCSdcg1j0OcUKZOD7dAq/9dEZNb0aBUUb8XmJyt+mG+JMDr3jGoYD/swW5GfBZpsK72aQRR
WqgQCfhoS3gLqCmB1i0sC0tJLVgw6EUULQxA8qLD3ttxJngg4T7iylPApRKns058mX9ylL5Hcnqf
xkazTyQ1SpymQuqHydKVHStSBvqBkl3QYSbiJNaVjyCXismbBA29mH7oBwTUkk5x4dMrYnWf667g
9VWYB9p90YbYlhWm4TIj9CkWjuOBYGDyFD6yKU82TNN7gpwSnln86QaBwFJFGebTpSNdWCe+hZDZ
qBMCxwKOHTuAJFLYAUdL43xD87h4X87lWoxvNhW0/P0is69825eG6FMKshVZfYssqxp7ZbB07cOk
MtG9LMamq48wuVTJRI0cB8DIi1gtaKKrfK5WuppoesqvRljONu9sSnkzS0f3M6e0jmd1MhEDLs81
qne+WaPxIOVDRu+1kIPdh4Uz2B/4kEEgrMFy3nMup9WpTp55eVSaCvFYqDf2RYfIv3mXVQGL8LmW
D5+ZIObyEfYt2e5HBS2qXzZ9WbPbm3r0Rv/2FlYlj+87AzuBNdcNVlKwkfZ1Lrko5tANKrk2WTqD
3ItS4dNSG6bMPlF92OEiotA8g6iFnnu+tyCtB5RI1wO7PeeluoTbrOTUCzptxnQsWYhPn8VpT4nw
XdxMSadvsgpfv2iCcG43WFONum6iK2K52MnTBicXavW5RmxsWv24sb6PRirE1juLHaJCi/CYcvhi
E7zAOqesB705F4bF4OBHmf70fvncFBpNxKm2w0vxJ7dfcEUNt5UOKtcRURBqad81u7xKCW1pG5yG
DStPZhyzQiPW0HNNwcqaxNO16xKQnN6geEIHbS/c/PKQrS2cqIkGreUsnaISKLa6IMS9XrTGow/v
AiH3ZlVuD+0jVfC2C3Zbl0LO0Af2NPZip6JQT1MedVskRg49G+yxCO7bu53hi2pxzJWTXNbsbtUk
NOUh2GiV6ocQTcarxVPkyB5zk/3AuZTVAjEIhde+t3ONcYcIZsBSYiGKu4yP8SzxlbgppNL31TpJ
U1wb63FRabz30xFK7ahSs+zG/hnTSwjaiCvQ/3OLSqRuo09j2U9NaTx+PVm98hnJ3t8l2ba9EDrQ
4/sxGmv4+Zs+CMGB5ev90f3eNplHeOVEXZsy9Y2aMeGAhXd9AVARv4C1ZFxb5CCAV/Rkbfhwx3Df
W+ZO5gLeDpFDfw/s50FQtiZNhME0a2L3WGWZafwPO7ps2pTjqsXulrqKEMK+HeKAaILELKckIh0C
MVjYJOK1qxbPiegl9gu+f5kNYLVSHnT1XwBt61ISexVoea5B9j1yMgjcWGqRNr5lt6Vz6Y2+Dn/s
ouJ4uczqiwbdostyG66OHjz2GiwfYYfaI67lP/sodgaKvitMl3zFwhZnpdyis+BIx9V68DFnyHne
gxhAXa/kZZ0HNQenew10aE397AjcXkyAaVY19N0NdhYlGOM91dJPXZaPSEbOYf29rjy4wB7PhErV
O//435TooatIdjirc8LKqI8NgG0U/3BL+18jAUiVMFZKhTAqISYCvOFFrizcMRSTseCTBJ9p9D3v
ptfkeVQyZSh7q712PT3Yr9b8ZMPWwU1L/DADWubCo+As9LeXbOXPzYRujY0qXCLtO7kZ9p1a4Pjr
knQmygSwnP24a1QsCOvNGnfA/djBieLDWmJvEH/eWr7DJjAHiIgpL1h/q0nVxsKTQs931NWMgpvP
Xj/GmlpUFciWwrEziCxt14ukF+HIaNgjtrUFFkOjSrIFMv3SY+iG7m1evEDOgnNRWzcKSDLhmagk
WZoI/nC/aObMqPoJ4Y8UmZmTAXaANtENACHvboBJFviVYI7Jqka6O6UtHFFELMNYiJAWEQOZT0/I
LYco+yOhjzlmLg9MZtaCTFQMZLsAMzfmexLbhoxXbSYmk2eU0mYJQhqf5JhdkFe0MerUZ7FmA933
TuRdzAynxkGXVjLVFzAHEOf6Os3YOgMYZETmSvBQSEKqkJEaeKbmJ9W2Rny7lpqjxCP1b45Kx4A1
Oxz8QltE5TWdkaD3t6qGHy9Sb5oXPZnZbeJ+9Wya+DMwDLc8TG0A25rJmxNp+7G4ec+CwbPTqFix
qHAbGcrhysoLwkQL/lzU+HgzIACiGurArQO2f/9sx7A+c2aZxcxPK/onpE00MOVyklwQXw5XbTMQ
HkouYdCu0iLL5gcNhioSeR0npUn9OULKvqtdooKiYh4EyJLFE9dGVosOi+zZouMt9Ypn7pT0JMjs
ZoSD6uMmjZDFSdG08CenRAQ/EJeQDSvarYN8o6JIXJbRf/VRoO7StGs02BIXGvkK+5eG+k7QkbcX
5fyGXZV/o+VRbXSwAq5Og6E/qV1KqHUzsvQWekL+U2v8GjuiuNyMe66Hw0usa3gUkIOwFzfsb/W7
nS4KWy3LKMQ/2BBLra2yQCawuNzSVfOW/xHOtC1Z84Aqn/rJgUhvkzXBDrWWnxllAJTqa4jOM4vx
w2+TYFiM+Q==
`protect end_protected
