// Copyright (C) 2016 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1
// ALTERA_TIMESTAMP:Tue Oct 25 01:51:03 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
EZClAtpno21lM4g5+EGOG1aLd5WvGBNE+9LppQNGdf2rXrrOW1ig5umlGTeNBeKr
KsU0PWRYYQpe8tIZKzKZ/ZXvm3n1aRbENC95F+SC2uk+g61bs3ITGTuAe189rzfN
5zrvj/i6tvdVZ89RZKiqRCa1lEUuCF+ppk85wDCCGDQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 25120)
IvFGIGpWL6xLeyGIaKGPLjAW7RzzIcwsBfx0jrTrKZHMahFvG7ORmCIUuNuI5h6a
7HfsIHP1AKCYU8qCuaDazLd3XVd8qGdMV2FdV7IsBEvM/HP/XoQiOUxqjEBqQ3wp
7H9Fpu700qxS9IF1pXEJH3eZ1CtC+qIf/QaNQqsChZm/7AnkzznQmJi7RwnD/Lsu
ePS4kj94y8SgavVNAZh8hHbKzqi7xfScM9fFYiP0DzyecKbcKix5Cx/fp9q7wBhK
vqKE3snPfsML2kLVdN8kEyq+JaRyKYVzU/XTe3YZfvsEZoDLz70gU9BWtcMAnZoV
Z9cU16Pw/MSwDQysjG2IPUsmtnSpf17gOjcvGCZA57e+rkCnckdHFoDYw9kN7AzY
WE76nz+73rcXCWlhnPW0cb+KqKltLyMThRp2/7zd1ekDhDGmaJU+yuFoGc1j2kGn
/bpCAeDWWsrqzcSOEKpNGh+r9a0Erxv3zApeOS7QsFDhqTVr2Qhxt1hySNgAhOF/
l7pRv/vodcodZRwNMyGoeBJeLhI+RKyng5NdUlyhBrwDDEvQOPF0WwxPbKF1Dt+T
qKrirkywS+OnYKGv99bdi+OT1MdarVHKFytvGyL+wV8NGUCyeJONSiKg55LSDORr
ukQGk4GcLxYVb6L2yuwvWRsNbcdYyNRhRePojuwxhcjWYJwm0LaX/AREp60mKx5D
wtL2Y1pYpuGlVBYIwrv50q6wZY1PUjV9eStzMM6iEMUwtyY9qpnwux0/w/NaWQ06
KqMYfdKLNXX34rIGrabDBy3hFVqicUVnxH5VbMSQ9YrQ2aMl3Ix5sLGUvM0OlStU
E3K1aHjpdmXMBpnVFnZGPgJ3RTZ5hUyEqCuheEWiOrwQkNEb0gwyxCnlAUg/Z9PZ
rdxbGMU1ZNldZN2VaMoT85BXddwIOpZ0CRL1lwG9f/9F6CQzLzbMprN/7BCRt6BO
r/7TZUxq9CRW9SZ4KnYOfL9aSMoExgQkz5u5OZHGVXDBi5HaDHMkixsMc1jyQnHJ
QEiEdwY4Yy/k9A+WYKkdryR/7MeRosd6a+KhKYgsM4/bsGzbzXpf9Wj32xYKtjqo
qpXdRlO+ivUWaxvIO57xYXDlEde72HVcZOKWeFIvkVqiGi+G9FwEPkHIVo3mQAHR
v5W4fAY7mr6bLbU3+EckMwXfvUPqBsNGfPwl+MLYCZv1Dgytw1bB5A8wONmJJX5m
nr391Um9gzM+F3R9aFojM5N3yAWGzZ8kEabEnd5jA/Z7rCH/4nFb64aHOPiMhxKk
qy+m5cB67NoqJrqYSemaXA3p09gxDxO6HabWPdWBVIq5VCGQZPdmt/L0g9uD+U1a
I1bPpODaGepdt3EAW6f8bfIPhCULhJAmGNnXuJZL/Olfz3/OUBGfVDRyumzEuCMF
il99HhjFX9Xh6CJ/cnvtjDSbMUBF47wbOWOo5S8+fbuZh8k5tJ9VS2oiEPQh7XA+
//B27Rtf3/o7vTkJhu/3UK2OT+Rn9Xqvx12LPhMACISXLMgaEHE0swQxLZ8Ox9J2
IvSXBHfrPLBE2X2pYB9Wc/Bu9/SJ5SjnQ+A/C6bNh+8TLm4n4nGA05ksilVpCBb8
EzvUnnEb84SlcZewk4aIKp5llLulU1KFmbYa1Ew8oMXySUI9uvhH9HaoN0+wLUDj
n3Omalb2DT0HwPlPpT6wrk8HZLIMRy9X3UWMk15zvej8HpuXSOinzhDPBFNS4p96
JpaSNZi60L2YPCt0STbAMhStPQiRYBVf7sg/jWfpX7HvTGU5W2pvTtirfuHyTQ4C
SNI/lG5PZdVN+p5xbGTXvNkSTu3VPbrrtVlyFMDBWA8cuJh6pnJn9OOD1qfL16KV
94WKWv6Cf3IndI9QeWXGwDMVxr1THWjgLOw7UFNmyduTlCP0glnrjMYatf/SyWSb
J6cO3rq6NAVEtKRseNcDhhGkKACLIqCvRFR8xYg80asrOKY2Ko+AX2582NCBP4i2
A4aBKPe6t4PHLPIarROLt7YnJENlaAlBRFG/TwF8tMupZlzjP+yJUqv7JA+8tp5r
nTRowy+F9h3P6tnPk+ZMYTiVXC2eXji1GWdDSfGqDj/itZtYi2/6P7DORDjDK7rE
0kay4QebaQgKrn5GXSK7jHCzv9ANQsmJS15KDQxgEQBuFVfNXpbzXiddiiQLn/tX
sEgOtHOeJmyEwRDfTIGhT6ItT5nwEQBE2JMW8MHEP9zk3jk6lefrqnNJ35+jdkPP
yMEhhg2PJ+SVBLDj5yjP5C8JZff2tl8meOEEUWmJGDyQaEl+nDHqU/5Al6x1IWoL
aUyJqZ7iZLGMNKs57TN6P+EHBl2Ermo/fwVC61wxHRQ5cG5PMBqFhDeGHlZf0jT7
PqJt+1CweyyGV6G+ecqSgL0sKUNMcisaj0LeYu2P22eh5HK1shLezD3BKLGDbZtd
t3U+WGwButwvlkPJDp7F4+Y+1oixezWdLPHU4PrJx4Vk/5cKFoWHrW844xrEgBkR
CN4SFSTD8XAeN6sao6lGoe22uVuoQidqHnjmBsL8l8twtSi8vhR99Zb37VaJH+Av
IICXthxW+/+2+ziuwvn+jyM+jV/j8/atC/J7Tfa5UcsOj4cV27iM07HHP/Kb4auN
5fh8WOwtk69DloNOxd9nekI1rG2ZL35NeGQ9ZL5XTYQwYTRFrlgIM4YgISibLSSx
uD/y8xpgJ3wAKRkO/qAjRJxXagfsOqEobalHHHUuWOb9h8P272ssO1bz23ZBmprN
iI3xrFWtfYYe/tn67UcqXL6PKx9KJzTk/hoCIwZ8QMH1AzIIgd0UdOhuZMDQ4u00
llMaUrZkD3ypZHTxvUYt+H8Lo6a8mVWs1vXQCwNAKXAL3dbEc090BH6VDNWZPhgZ
eoxrWNfrKsFtDSw1W3NiUloVoTjgVHOtpUdxNtmdu5CK/h8OiIkzJrMFABgmXayE
cyiXTjB5Qeb9PqZyyP4301zx1dV/SVyDW7Vy1kZQ2WTV5MAHH2c8fyQ0sEH1W4h2
hMhUY+JCNakkKRF1Tehof4mCR54D0aeJV0NHJKbbHCbsIppUMErFv9zLkfyh1lHZ
Y4064jY9Bf97O0BcLgm/Tjaf30EsVWTfCsxayYBHgIpYT0SS3BLf59XTgFWU60tx
iS99qho5+AjbAyS03V+GIY95c8VXgby8+cG0TrItmq3Aigek+ZdStwBoFkdW281V
SLM5m//Annh3pEc952sCMtFdIYeIGGAV/CD6VIH1c4RD6v0AiNp244lzzHv44q7z
+pAgdfpq1RleJA+dqxSkc80YNyFfsdEDvf4Zy+t3OOol1atXtrrYv5rNlb5eyRiJ
8OhbarMdBy/uJb4RrfB2KNj14imT1Yx2vZCuXURXk1gokG9bvBDm9fsBRGufryUV
UdntF4SlDWit0zhuC/hG6jaDccV2ePiPflKUHwdYnJSuMJf2hE7AYS7pNocrqZ9S
IG2of60YVqupKXqPaescZNOGBvL5eKfBxxsv82B7JlRo3+Pr0t5llbmGfQ2u7J6T
i5lvm4h7x7FXPxQsanBYjlqMZxv2w2mZYAMRbB3qaXwtPAZxsOddyFA/psXyEx44
BBTIarvRO6EEZ4VAAp7cYuYDQ+VaPtWbLy0tW+u2f46dJiT1FRK2p2v+sdXB8HFJ
S39a52QtrUNeqe5OVtOPKQV79dhJ5lq3edPj1Ot2R2NGacpqMa6TeYfMAmuuqudX
p3kh82OX3BcKkN6tuqy0KRjQhf5OXcRr9MhsurP4yfM0LzG5a4s+eKGz0TdkMn4R
7AlispCm+GxEDtZ4WKh4AzgTSWfKSVnKuryAgJzIiyOQ4oraOyJFJ+jU/SPtIk2X
Abl3Y5+J8evBCwYMA1vAYmEYx9BDXgSvpDIZGqrPwtmif2ZfCUJ3EkhovEQ7NqX/
RaII+ddT1RRDKy1RpNdSQaw2glway5UipwQ3cSzki98rX8/Td99aw/Erd7Spdqws
Zu9XUfep/A0ZbYjfnDdDkex+8jMSqDu5StkhZbJT6trd7fMxN6PCPBLsmHGWCVfq
wlZVYREwJ5Es5dQ5f4edm9xixgOKIafcyxeDcI5lyjRGHpFTBGG1tnIdBL1y1mOg
MgjgRkJqztOAp0YOtK0MwPLDlpURulZ4uMSt13LPs9d3PZD+NdgOz8DPVLfEQNUJ
fn4qWzCSXzJ/z/xRechHjvDnUix6vCoMXeiD2SXPyaOQXqQoGWZ8iKUpJrA7gPjZ
tC4dPXaUgonwOX3jlhCBAw3F0EcvC2Ln3zEvIkiOiSGB1jEMlGR+De76g1/SSnaN
Jg/WiKdGffIrMsLSp7Ipa2e1Wj5iYm6QIc9GpE2jCEyzy87Ps4mr+geOxH1SdNFT
haL61NBHKen/B+FOsiW7LsTRv2tup5bU0qIloPHfFgz2cnFb7Vk2yyM3iHQZIwBo
XtKddpkZXLLwg21PtvvwcyZyZdBRQVweFTuGs2YddtnOL5rZkxXQ+jRQCBIlyc4G
eClHLSGPiBmY2/lLO2HnjQtFco0RSi8vGlVKVv9b3VFLYe5G9eWBWaHiF0/xMkPX
HtzV98Wp+HsjjCi8rd9esT8Qig4I4X7HGvqFLDs3pM+R9GT2bRLbyE+r/8ZW3Ok1
g09Q2NFORGB8WBHpGmSrJ7q29q21KoGXVZVV2TNqeKBXIKems9W0AO7TSZNeaAxB
q0kZVkq/+YwleA4kpZZmD9cnhjBv4YJmrdP8DpVGuS4wVF87ZOYy6Z03Qjx5eODg
sYJJm/JSsaVHcbsctKu9fe8u8iWlGaW+EiOl7sUVDOUEoPIuSwSUQzo6vgOqcdRn
hZqx+8WjVtkfGM2qTPoRGlkTr5k2qf14nsPIVeyAa282hL20CBN2SeDLHZ0HgP+0
fKrcJ6J+D9DNJs6qwlo2VWouPhxaZwp7tw2cofMS5se06MFx2JO55/UQqQyXRgZR
mPqrtM4qQnRm7T49Ey6WUL/bZltu205mXP2D8tR17hcyJmTijaG2kxQ9Kc3CAtjB
hr8/jB7xvR72KBRcBPkHoX0u818SpgTQnSMmr9gC8neMla1sSc1qLiUldrgtDjYg
0laFnjNPt4qoPlUrCxoXlZ0OUsVF5r2VleGkNRnQmahbqgQFeTuxMcjhqCT3vIDa
VBhFUwngF/UmNb8GhM2jr/pt4PynQcsLuKeeL7AYUDbqXvS0KPIr8bnHg/kSh6XE
x6xVhkvcXaXkOw7JzbqZ/DIcXCl/kkGJ2pitJdBhpKZuF5RacnvKSf8z6u1vfhmk
wZSz9w3CnK7FX+pDigJFbO0bB2Ip2WHLC6U95+WN2vDvxQfEhW1cd37UtirakVhD
iFeGno+I0oNAO5shOzAAGVRyMf9gTMz/GxneV2lV1MOIjawwCK2vsNvX4seHypyY
JWwRpkU/6mx2HcsFt0vgmy8+ZrT83oyzbagiXLVQXhRtEjE8EiaA2CbdfqTjdgxI
UrB6+F4hGA5nBHOBxMi+VGmBR8dOP6LTME2/dx5i3YQtoI8KR49xHDE8ovotugM7
tI2WYEF+37qn7eBzjEraqvJOi7cJMbO89zZq5sYk5DuigX6QtfsmMh6wwQuLZq5v
LHnCoF5MINubGzeAWsWnIQkR6JvFrB12d3OdVEcJ7GCZHvh8YKorOPBj/4zmF3fR
QKQujTRNEinB23j5Iyz+QDbch/7KGqoiqB0bhln4n7tZ+6jue6Ktdrw3AG8Xs/FF
jh+YvFiwWaoLDAW0eaaAatoc85KtYAmVW+RsOBrF091YQtKZWFt679Mu+zaTXTxw
7Yy+kdP1s4L7U4upyFkltrcGM3wZI6sw4PqFR+PC8OM4r7TDUjnn9qW3/iFyU9cl
WWI/zbLDNbXK9b0YChzEsPlsbA2xilBn/nsPypYL80o7uLmOtdxBEjrRnmnXZnOY
+Mo+OnOMsL1KWgEaFVp4I68NDc6NiSpHUGdoTJ8k3481EMqOD2+tLOBoBZcW8O23
e8bj23TBpMaUtK+uxBMpW5eURAjEw+useahMQ2Af42W7JRMuXwguHLJCrHEpo0NI
sApzjKglHwFCsEH3DmvDUl3JKS0DjYPl674tvA159sEdlNJIemj0Sp2f8MZaROde
5VKXR3UDTLbmY3ycT/ose/z0KzpmdlYO8rPW9CK7TRsGH8cOuEncFl4ywBq4t5Jp
3CifF5IkpUOFaLK1gk7xvlAw4T3x9Sf1XjIRXXAEzjVeBwGiD4K6xhjyUhvEO0+Q
Of8G9REkvqHC6qvltEetYL83bPEMbZFBqnZmvRzAVPYzE4dwa0H6kgGm7p1yciZV
mwlf4Yd7PRAPmZ64ERHdqSWc+PaQc50JLsiT6Mpb13MYzLiwfwp9Wvbd44qgMR2n
dpRjs67G/+LIJgjkdzVOYxUigPGYSMugpC3kM7QrNHJi99w2rBt8ce61q0IKAEBt
erMSkWdj+I0IDt2LfQTn9Q0M4IgYSCdBdNCsVsMxG5ItHEZbfabLeUGRuKW6IQ02
pdCkT+ZfeYd8B6RszAHPBw+hwALK71f7knmM0LWN84R/NrwDX2xg90TMUt9z9eQa
ytT1aWLCfFUbc34Xl5Ea5whWy7TSGTGBdaHfnfDKU5NJ1TU/9F7GhsafcMwRHjHu
VvEao8bYzDX3eOBmjSfIdZrV8cl2Di35qsdE/TYoLJF4tVf1dEWEjCwq5U/jCrk8
s8KKMxrY/npV8WzHTA/H0SiAt3AECsyek/Ke59KwxL9dU0wd9HBctuc56C7EdyhY
5wAXnCiy7q63AZ55BFdj/Jpv/At7Z4a617ZuA+mGGq/Tu9gFDBfSvrgAR/QexztK
npZf5l7RbtAQU7n/13/mkksjR0rDW9zc5fUUUq1rFpPAdbfhGTc+yz1NNSoVyOSF
sSAJtpLG7eNfvsu9JmwOweM1kGNkXxguBi5poDpm083tYgZaYlhh4gThbbnzVWiZ
NpmaAArDX8HM3pnj1xAUD/yuWNPG0DO7FOplY4Htnal6keteW7AL7ZrFzX2ZaWJF
eEkGMF+xgqEX6AyAOAT8KIhXbofrRDmFT9GIS/fTk2bxebENO95xyzT2j+GTEEDO
PDloK3VwPOXE2ST+BAbzPQ54/xZWQpFSn3oJk1mRL//mUJSqKbJmG7WZxPv3WOYV
P9AtgcuiSYGjd2oDhJxTnaf2kNyGUzkmMJeobs6GrqmHBOP18ik3WkU9PvSp4IJA
JDqDDPBPMDUn/2Z7hhgVNJf5MkbjTjdtnnY8F431Ze4ZwmU/esNhFRbEzFtaQ9JA
gi9o7Tj+u4r/BuwL2uPk7KaBahusUkkwElwcMZM0oUUCf3+uFi+jYMRLV/zA7kd9
IvSl1+fKvk45gvWP15uvihtPFhhjGrJy4lAUQOmFytk2tN9dImpiHgKHFsfDaPTC
v0wEOXFnAMF8QCeayjG4adWBkySL8s/GgWOtVMgJhYhbdymlbHrqwiRIZuq7iGM/
wVTWUpeDNlr13XZSyRopggvFxG9UyqDsAbb0E4pUInCF66PRnHIm0L50u+NpykBf
1XGUNCLVudrEGdg8EvBW74hjX/mfnOUCA8B/45sQIfOcA59H77mbHlOLvpv3dVzD
Xsh6MDLwrNSvIwg3NqhCsB5SqlNd6sGOYOSOgV1eafnYjGZoazkPHIVeRlDX6K3p
VXmUcecL3MrGS8JPcUClh/Sso+xuZFEu+8pl3tMh3Z6HT0a87JAVjDZet2Jn+1Q+
lY9huNwnVaiZhGyeL4HHNu74yJ5ex2TzM3dHHGWE3ngKrpC20IB0rd7B9r99URdB
mCfy5caj8l51pwEoS7f+IUxDS+oKqOAj12XwsJuPf3ffBOoezBrhzdkQRgQf0GWx
MZy9zua6+nO+S8tf24I9sUwUf/lQr5dJR8xU9050nDvcVkMWFCzYN6tMx6MfmOtw
PN7J0nQWenEpa6UojotVht3KVxw5ffKwW8ICoZQ1m/45aRJbAHqfXkSNcl49S4h5
u+jf8SsXt11vOuybKeeEUzsj6jgb+r4wLm8o4GeM10gZ72YHdmmFIuckhcH2WldH
wr7tQ1zyKEFVepwPUgx/7J8vLzK372b8tKWRjBkPak+eRLSY2qYxYDQc+eGp9+Kr
6hp+iUxNR+znQL7eFGbKv0UvYJX+fKChsrbAoc4HYFee5YasejMOAfL3ob0HJAd+
6yZsSlDLt+bWwBDGuxFLwVEpzWvj13LFyivW1bNNwAeT+Ew/FFyXQpXx9bktwf0G
tTNVIjy8g/39PfS3t6oOzS+Gofi93KTM54Y3wnR1jFIlj0UZGQz8ammjgcF73kLC
ehHG9LjOGQ0uSGKhstTR/pbQFuhTX3awx/IBsvkKzjQF+WStjwd7iffGXhC3Ru9A
gKPKPsNcWkcFqe/CbhOj0ABB80NnrJc3A8KQ3tNzn58BFGgiqK706vo0ZwOTJVyh
QSIy03q8iLhTBHoE3Og0M0jx/ABVZ7CIEDVFXTPH/ULbjrahzxKVCuJs223WoNlu
xlmYL8ATxS6KcIVoWZLMrzGI4InDoEl/AAprHMwMS6VwFkrWeOnimVpaXfPxNOWV
RSi3lvAEdRw5v6O3/4PhWlnJWO7fg5bOwseRAB5Jalypb7QN0JvHclOt1JBkbN8h
Lf/K6GM32o2p4A/hZHy3mJeR2R+7ztQIzf4wETaGZirGHXMwQLYUimJsd+M8AUS5
VhVn1bv/eC5/Npz/BaMltszTbIF8jOBzifQRLNmxG+pH3cDIX2BJJMkSD5Wbd7ga
kR2TJmjSMvcfAUWnFQMrT6/ZTZXNiZ5nQ0nS3cxZJ+DaimFvw6KhA6WZ/sghnIPR
bsxY+ZZMwrBRAWVwmauEvxP1zneAlEJquCUkkbn2J5g/K82/dxH5hFGml75Ua8tX
SV12YKolPCxqaEti46ZZi/NHtnOnckiIOf2NLTMQZKcjo/Ol6wRlcqj6u1vIVRPe
DJi/beTfoxSNiDu7NwrD8GOmlU3I13paQFp0WyNiJfY8gm7cHTZVdPYVl6mRaH/B
SvLJKfXIXWkq1l9PLxSu5V9Tg6HgWYSqxxyHMDrOVB2t87VkSRta/9dLTAN8swYq
+izAgYs4ulh0amXdZvRneZ4Rrqn/cIjt7jVc+x+hsjfIdgAWos9pMWWPLl63AX6X
ouTxaeVxShXdphCOeYQ9vnxvAvnTviN9XihCKe0NTgQ69AGDsuCb2EfcjMmSPCsT
IMx+aJG42d7UJ/pIkaHY05UxwN0y0ztcnm7dcHN552ez8syuexVCzYuMT+SHcIZ0
CR1HMEPCbWy0oMnZVSQfPh6ppY4oht/6O7MYPBbSm1HrceSfZEgv0R+yfZG5jCzg
vnqe/STw6trtsqAxpaiR2ZsHe6Gfs2umJGeYE1QmwaPyKWs3rD26x0m72/Rb2oAw
cA0gWctKhQYSOKYHXBKyv1ytPcspNfWb756Odh3w/4fan+96SjLIcGXGUCJbFAfw
ClfJhpqoJVodDOL41Ntrfs46B0KQOKSFKQVHkyOP5RREdWZFuzwrlwjpeo85ib51
QnA7/bcWsfnqbA4BTAtbtt6AJHOnol1xUH8ud3U6hy1QkKwYWlv7iPGFX9Wf5AyT
agbOKU1z6uqBmtG3Mo3PZD1rAgrqDM8tj2cISo+8gxIG8juhyG4f7l5AbpsBrogg
95T++yZfHCku/NjvU5NkWhVpzYFK1W52w4huYUvRYsRYKrBa6von2j48IbC2+R1N
gZUCU3a1mxCyXI1iOW5OZTSfImA74tjpGLp2XBZFaYVusnIexCCfAXOSWJNPJFl6
n13DQA81or/tvQ4m7SZHPQEq1x3EGGbbREVZp4yFH/fCOqpNYSdWpURFoj5x79EQ
HqS6TozidgWLA4usxp4HpsDy7R8aw3EG/BZbzFKevHSVQc8/xZwPLTpYTqJQmW7o
dAaT65t7pkMOhYCofX/JAOHofvNFwpomSCnG2dCxs0T/Bb47M/lMi8LPmtfkgtMJ
6Ek7+3w1FBNT7KAqzrj9iEHNEI/I73zUseKVwRs8f8iJOhlcaIwFgPwwEqw09Qog
bvp8o/623V3CVxjaNEzkJx4Gl2VlW8Yl/0ddyeQF6+STVsLrc1z4JTcZtCr/ufsm
9N6ignFJO7fSEPCfyeu/ZUTotRJTpQODpMIa+xc9rgbrdNmngrh8b6l9JqTzcxXo
S39pdok3QWlDHO7nBzjexQMVnaVYkfcX5aNMdpOZf1fFdCXGsWlbPfsr5pCXty00
fhaRluyq1EIZlmzR9+o0cexF8xKLkXigPw/Nqd3yiKjZ7DNGlHRbJmRnQoOBeMn9
E5Kq4sKD6+VGnkUvSVGdr4XI/eaMpQRBh3RgeXyVRZTJYtJnRy3f7iJJswCKeZUE
k3YrwHw/ZmoPFXoLCpQ/0gtXL1lKadwXu2cTRxdsyhi8PHiQ/ui6n8c1WdstlTXL
GOzGnVlZ+c9T7yDVoOUAI5RUsB7Wku5DQSh9kTiuNfjIJe0DA9HK5PL9IvTSzEKk
lX0g2uCqm/a49XMFgIOAMd+rMHokMRhFywtSRk6K5CrLLsrRF0aEkahNXkLY7jaF
M0PImZZN9lcUvaiVGN/HdninFc8jyz+cFQrv6UIYncPNhC7QgF4NaD6MOYaqUyZr
Vb3pvkQE+q+qtECXCdvfNMqeP31gcPEGVczgbKgtZHPMAeUqKFGK6JdnsfSONeLB
x4BFp8Gfjg4Kf1xKvVy7E5nqxGw7g35XKAVAB5vJJiJkFMncgLowcmV8Q2P5/663
vI/dUcjxBG8TBznt46bySo3djTB0m2rCTECxU+zSsxruSTNK5K+TC3NC8htpUXO0
ppmyay5aY8DhiYNMFUi4Z6Oubl/w8g9a3j6N1e1eXykkHCmc7LFekMPeuX+cWSsT
VgciHQdVnf3k5i0Yk+Ulf0S/vcS1wq1CxPfDY49IYHtgrND/7jC5qAdeZjvbKDlP
5IqnyYfqXNEJGNyxwqEJPO/yQjwJASN3F1QwwUGQqIYMq0CH4fbkKIbJNUtglPMS
4AxSZTwCyAxNCVd7lWxg8d+sEyxs4+OAhoTH2pyVRKoZfXKrAedacqXnJg16wtYn
qd8cO2msmUuJWieimE1IWftcxjK/zzH+iXtQHlH53hIaRGfELGl2MKMvBCPweStn
aAyEHU81B1sEap2UzBNQsMeDITrKvcjdebq43DjoTtdKFpc8NsCfuBtsTFPDdwr2
9pV2kKuB/rQuMdfa1jtq6KD1/dH3oqDgmXKPjWKMvQH8evWyRcoJ/sGYpeAYmg+D
kjbSUasndFhWXgzaY94o/BukbtmO6MBEIdhnb1ypZqD3HUGy8rcasLPRFkSj9eop
Fce5oqBazthtohcHAvDwB1HM7B84HOvXBe7AXlcPwwRpl3+fhjgf/OK242TR391b
GbdMB8Z8YgflsLwj2sEkb3nzwjDc9x9S9QnVwgkD74abh67AS4DEeuxPqMufOMfD
Er9VQG/AhwGBB4P6bzlW4T9W+VA6sMywHzArBxeohF3f0Kb0iWjXwGsg0x94F15G
r7CuUUXYnbUfoVhHV7dGgDfYa5it5oB4W6ps01EX5YCatKONygPmNr4fc5TJsQHK
CUj+/XkVi9PvfH9Nn8HoEca+HkOQLlR70W+znn5Ns9fqQm25nvkemMW50EX9nB7j
Uznm60pLhoj7K2puQxjCqnDdNEzrHz6mDRXnHUKF/VGSEQASMUToQAst9OFRpFFn
K4EaGpI04NTThxfTcmxrhDWE6ajYRNpNDGsmqAjGvEikJHx5YnkoURHpERgesu/2
MqunXpLYntT60YCxqFr0mp9ziu2n/O8IJWyWg85p/k3ltIwV28k0PS5qCMo6Yzgb
5EhefBzIZ/SRgwOPXbDU6PVzVHTB3vHCfxN8EkQBQMV/I/7PCyLvudFXqs0fqQVb
fZXb67MPYAqkQop/BcHCdP1Cewo7nJSNVKTTdzhWbcKF8z1zSrYyHvh1pSvf22/+
oC0oOWxlyKY1D5NyRWOPWdBveJMRlYDoK7fWgp8ZNmlu+uJhQiS4PE3/E86mqZfu
KC5kK2E9AiR9LfIqsUiSWnIameCM1WeCGawhlpp/S6wlo77d8qs/WYTi3WOPU6H1
w9gzTlRxyzMWR+acL9jzuwOLvn2UQnYlMerRwqAmV9sm5JYBf+YkuTvCyUpxPImX
cI9MRoX6zxUxCuJcTX12gxVMi1BfPyWuVL/DVJBAQw9EGg3mnXrSSlgzekub0nAR
2PM2RwgIDT5okCtLPVcCkmrtq+PqD+bgPMDOJ14+gD788JL4Ev0qmLL3b4DpfUly
cBQ0rtFsxhl7tURRWiVBSkYGlMDzXuu5uxRhBeD8rzTrWh7BIyBTanfbj5sqJltN
VYSMNufpg8XlvViWf9WWEiZR/27DxuctwENZicg7QBgpZM456tYC3CEZo2YlgGLz
XCm/N+pU0WfkZXRuEsA7IfYXHJVKGAScqK6KJ/l9k1VuSKwHYsTP6I+zof7sNk5r
G3JMDQg4lplXpuzcjeEoelNykH0QqLDVvA0uZvs8SkAGV+kJfgzNburkSEI+tXk6
9h+8h5ITMEL+jO54WS1TaZRoWwBOvN3O3Xp20zoBWJKm7bk7C9E7rxnb6vxYr1YJ
5wPqYQ21XB5BtbwmGTd1qkMvPTRu274en0FvtfMneYRIqiogFzdNdVRnM5punmcb
KsnYu3PoAkHcAIkY8A1F7IXcb9dHhDi1yPJnbCbsCcwcrsDwnUCywhwJ4LgeQOkF
ZmCDQMhZ2EHqIApF5uezlF8dHta09QHENRjvh1EZfDbqOj6bkZRBgnZU7cGp8tLi
9EViQXFiZVUH4nSV4m0LevLpdeyzZs33BE6Kn+c1I+KovL2fTi80+/Cf6u83Y3WS
Jify4QK/YGwKCIRq5NuBpx/qoEQC0j8pUvVVQD8F1iR5q/rQgf24innOuSJoGFPK
2E3MkvTsWHw21N43U9oyh8GgPg6atPafZJHESNRSYc/JECXvodR88bE/JgvlmEJv
M+ZAro/nlXUHXy1EEyhwObVAe8h6X3zDHDhcZAF57juotGuA+rvl6QJeatpamFpL
5Ai+NzC14tE8qXUZS8Ytd6Ej7pWzLmdbmKrYdLDz97gEqVOhJQGMu5gH9JHh8V1D
SO8GHG62lqc1oP++O56BDCeYwObdHJriH3ldfWSvrLHB19ObGHMmQZnyc67sO2II
s0cXgMKqfFG9ZQrCpvuVPehSrrql44fAnl6BRROKNBu/Yvkv1t2RxaZ8NqCoXpbo
OaD1j5UuoLt26EsWkaxbnXrmq7wWh7VLZ/VOqDw0c+gzR4yL6v7KFdLxJj0zhsaE
N22Ykehjl2HZgSPjHIc9NN0sVJoXSxwYBvO2ekGj7USzdzf0LTYSFSvRoKNfZwB8
tJSgiCe3ONAz9hGWfq14QHYYSii07zsq104Xr67KH0OHOGqtEhECMTthsEvK+IBJ
m6dfk5zcyxLhcTCZbZV95YTJThoLZ/uRjVI3THCQqxr9tiAfTUGD3EyGSe/RenUa
pbjldIIkck3Ke2JkJ4IQKcdUBQp0zYPkPjNp9xsKD+Q3YtIpcrXiz0NpKFkbc7X3
j+8IxB+PviifOuYntyLoqr7hbb1unPBO1o6MNA9PLCb77X4SIGx4SRwqq+5IjjGe
cpsJXLx+Ygl5KGgXVHgqUbtG2YgD+70Qksv+2GL8Jpa/SQf70U33zDXULbzB4ww1
EhFrMaVIA1Btiwlav5vuV1hSr/ww4midE4C3XwbzlrI2XFbJuT0e5+M75hm87R8Y
fjNDL7EkOhYsR7RAG2NCiRekSQgTeJo22I1oX9F5oqOPTCUVSqjpqmnPL39O9TZk
32FvLzMPw47cnr3gG5xwYantINa0MuV5FUMZt9jS8K320RJiiGlFsu8vhGu1U4/h
erk8cgSbEwWhWUreEIx1Tn5sm3T0rZSCY3UBLH4v+p4VCIzavoIVRwlIiogw7jyp
gxTYiJJN4A37+89WZ/j4inmY+VmbKRR1U828xVt060vs3kPwT7M5BIMUCTLWop/9
4JdCHlyX3+FR2ijbOlDIgriypV7j9HyNmtjGHDbiK29BLs1xagciyJ5xShAV2LfU
0bJ17ZSfWU2k+PJEouYCBNk7BHgMnsLZNMuZX4ZvTkvbvXIOorsI2fFPp46GEK+I
DjSOsIAfQZqsQbS96WoGD5LL3K4XWWHn6wcdD2Z7pdc9eohKX3D1iaLBpGP3u28a
WF8F74plDOORkYyywpgkjSoO0UygJTyowwQPzd0YkVdw5T5qbZQzT9x9O0Hs4iZT
vZt8w5GJX7U8w/PAc2+8PrhLPhJUNsxtYhZcDZO369DnW8tnji6CvmC9A88rVl38
BE5H3Rv6uLqu3qz3OHjEahhYRYxm+ZAS9Jqc62QN0nw4YSTR8IQjrOZXWrtMLG5P
/WWuKXgY2zvibk9FD5ORfRhxiAd6Lvu9Ogpku0DG7vTfrCkh089FiFU+rdqHX829
zV39dq/vBOEjuJIiFdDkDP1VrxlioVAKJ6UgXeV3E+c1/5whambGEUHPpFZxjEbh
ZxNnOUBmfFl2550GtUE/4QfkNNmyq52S36RGR7+es1iQUbWy1w26iTwHZBfDoMVh
JOmGwb6xtium+Tc5yOIQvtX3SJjR4FvFuAgD9cIVfINDkb4x5Ayy83Jj1Kcy9naA
1GvHkmsfbIP8VFbeQYZke9kFDyZM4oFOHj/BeXGi3KfAfp6seaFP7qhdHkwqjXLp
P1oKidHUe5BD6oa5ElX55Uw4g+4mj/hM6Mim7tFOBpYJ13VGA/FMgQ0fQzuENyZZ
r2OQ8uyhrV6zKR6JPPDyygD23TZfS0MPjiqmaeGOa/lhunqFo/d3oF+tmwo3KrL2
HckDGgwfsu+sVoery07aKzKnZk72Wwme+qtQHEogHL91lq50FjuA4hjIPt+cWYO+
cYUJTnOsq/S4aBtLEjuYPShvqY5/E2L0DmopmZjORUA0uPT+DtX7fH5Ywo2SMdn7
wAlcYTCnhQYsM06gqeQmMxnZf5ysl3FoMkkdj8yegygdmcqKPUtPvSfDUDCvHvT/
c/Zi9NVjLd4mWtygq3AagCbtmiqU3Z5dhuuyiO3ItgQTl9ANy/9g9KxN1ii0mLwt
ubRYiDIcWzfSohZLUXEBtIW63l5H/waJdOYA4fVyVbIAoiBgCFoiTVRSe/5lOq4S
CqyBaKWLMKxsmOM/pqAMue9DV2e7ApLefasNxoy1EbgkzJEUqgfEGeeULKdD5JK6
mCnDkRnACgwxoShsjCGH+QceUNDk3NW/eDTVvVna1023ieBRLpxTxZzFK/RMErgY
VZ+6x9JaZADGWqBnkd2UatLs3+UPoY7kzHWv6+p6f9T75zQCyeDnahlVlwofsjAp
obJHf71a12ngD9ME81/KPKLc3rviPV2jwQ591rRT2SUqVHz41urz8l1lcDCLHU2Q
e+7o9vfKTWhCImmpOuRwTVwaMsmDIk5pVp3GElRMtuQmSnq5JbE//x69wwgXLHq2
0RiZxwAIMGyc+vQVeoiDKrtlf3R+4tZLqkIwcCFjxmkB9oNiUu+QZYdSbO3jQ64P
K5B7vl5NUOIk18akE2mAqL0QBGbDbXgxHJMnfsqpE8WeXdXFvABR1Ihm9lhPIoZw
IiH4sYuawehysjjPyvIDDS5t8Gkel8/cEeGK67Upz3aTBdJ14We05ROMGqJlsEw7
TF/xmlpR0YYza/cdMeI2zDVG75RDMKUpBsbGly8CB3mBc9MM6FsHWj1WJ6LAUKla
dQ/aSpN/tS7cFeJmd+7LSGr0H1G50HgIBRtNa+KUD9yOzESCqzx7/Ye8mvtNU524
lqhsb22qE9F4/5roRgejoBtPpKfs19kvkQPAH6quJe/0OgiLco41jMJuuYAFs1VR
aObkhzzIWvtF6KvgJtqLiFqRU35C8BcqfcAqLHPXpKhq2qcH6XWez4peQGVOYc/w
Vx+W1HJ45VyQjYwiDo9EVZrqpjmY7ezw/JLKuydUWu60g+J/5Q4E3+GUu/STIbmR
iOtr2NOZfIwpeTJsAp4hiux8gMKWdksZTuQg7OgAsJGlF3jcpjHiYPSslYRr/ZwF
bXuJ23QBOSN/CKTHZY0Ktl+nU6FvzfSM6bnt3vW/aWLnGZsNBaqFH+Jp4WflA5nN
8rrKgImfh9cK7AY5X53qvz4sUeCxXq7fb7ZzQBeJf8Mm2eGFjJl/Ht8QDgA4nHdc
euNBgDCCRleT6+Kj3Y4PtwUxpaRXrDqvy4rB1xxcR8ZwocX3y5u/nfZSwDpUUB5l
bTVUPOWyFhYN4oxrtDCY7vTAkXxZeM7i1zcdEfQ68kXX6VtNe3kxG+NDZ+++vVzy
jmQUqWAyFvCvSXUbnzCuZezWDUsgHVclC0YdnOPevxwrftFoWCCUQhVB69ZQfTji
Ob76F08zZcTTLVjQBFfvmzdPYUwtVgODTZy/aqVBN7TxFLN5M5u4QoDVv2Q7ivlp
MWn8ElR+ynJepyvP9sA7/KcIMtx+4gMYeZa149MP0xQEZc060MfrEDCDMIEH/UO+
lnX2Xa+RX4+JyOuxUmK9k/h8Q1zUkqDR/lfZlCww4ZNDY+Bs6DH8QP3//NP6GED1
B+ycNQADyY9b4At4V23S5VxmhMRxU/PedS3eslSUcnEfAbQXUAuSrzTEKWKuakgR
LRfzyI1gWTRXWG1kyDvZeJS/lB6htXiYJ6+bL38yaloEseRNKcmZf8qe0PnukrcV
rHtAuM7/FfQ/tSvCm/NPWtHkNBJJqM6GrVVw4vmhp26mSnwGh2e/Bgxq3ZLviTBL
gA8njM78mcHU0GaJKKxuTEiaSHK4gAribQj2uh8reHppD2uIx43R7x4RCu5P7uIu
PAlybuWC9Hbp4bxkbMFhTK4vl/n1N9rnNf1gGI3Cq6JsVWuL07eh7QKlaYD8Pefq
beqtG44ZeWCvTLA/DorfNSa4YM+QNJdJ/QA9ME2aNqU9E+mGaNmhR1DeN1aepFkG
O1UIKbx0KcKD5NRLJQWzzM0ZFsU/xmMEbNWWZ0ZYchsyphevvGnNELfnrqdd8lIa
Tm3wVNgZ/5tEHZ9HJxJuHSTPFyi/FvMY47kUeSI0OyLWQggPVz0RnOnngVrurwvU
/AfuwAqwPTPplExLwNb1QzHti8RCNS7vDU7u/ftuvP1sdTlNnz+14wzO74awkZLb
ff5/ADHI1mQnaqoAbQ+6b0MMXNZjNI9gjeneJRkfbdcSKsa92sDWyoc8IlcBW2EU
dmqwQVcpg5fvNQyyV5fHCwpdKtEMfbjfYBCQ8F2Xntdn2vrmWw21o9S93fA8R5Xy
5apNREN3E66a4McBmFw7R9gy1kaNAFhkPUy77qU/HBk6V8Pn3FvAtnn5JuyEnhiT
6kExvOVDvTCDtdJ6zllzUoOunjjtN/7Hp7PKSEs/5QB86vqBox3tZZ22CoZiv+9N
8n7RZ5NCl/3P/FG+mgmb0m2TMPjQ9j+47CGxwurwFGY0ksdUa3MgwtXqUypoeSLj
D3UwKmO+BSibk7Hf81a+ezKdsJSCX3O0tHLMbSnRSpkPo3yJIuM27iUecepsJZ7q
4OqeEW5i9DDsPDD8UpJuR5/dm0/ZnsIqFUhwtCk2DR8UXs3sOntJ8IsNIkkvr+vY
OC4rTEnAwzuwtGPiiGt61PQdooC6XWc2bm5s7hawv23Vf+OoJT8N4VT1oCugzvge
XO+yhXO7SuTqWUKsJ6GSu4i0eOx/G//Yq0+J0h2anVj91VFOQ3HS6rssz2FCdOV0
znH3usjFAH5YG0peBrFyxvP2ORuXQWEDMni12yF1ew9Hs03OXPCoTaR1rwP+94mL
OmQQA2VPU6+Nv9eUaZrCSBQPCGJCdseGFYDRj8eXqXJZsiZBLsO0MsQwMcIHOYvY
hxYlczH9CCsDVku4b61M6pYQyH0hJszIs2XzWIRyX1WAOn2LhNUstF3y4WnJ4QeN
p3SXxdb4ak6+DzeDtnAWcLmrAKgZ4ohe6gZxt5NvFaWqiVS74WHy/5OjKVM7oDVG
ElTIZIGI1RRgn2aqElg9YY0K0eSwCwCJ6P+tZz/pWHqTmHJboppetdRwvbYDIcK3
h6k66owVrbyQC6SnMPqdkUIEEOqwFPF1Z00fvivu0ZUe2e1IOqWIsqRNyZCLIzl2
cunniA9ihqL9TsTYbziXmWj/uDWE5D2pd68OWwtKDvkAxfmXrFw4DeR5Uo0S4qB8
ATM+ZBlUV6JAYqIyWxHoXgb1LS59WQ6N6WOqPI9E0wasQ85QNniILTFREoEpOxyK
+uMQ+X+vpgzgBv8R+nHoouKHwLCYHaZ5UoVLYkqqH57LoPdOGovXOUKC1NLou7mW
jmUNcGJ0Endf9fmXO9mTeurb5AyXpadrN7aBcHfE0sIdk7BgYClKvxcFTIUhDrUL
dsqnbn0uaQx57M27DNl3CS7fF3SeoRlET6saFaKO4Cwn4m0BLqdYg39jgt+SChyF
tUgkNZXm8+u2NqopozP0UX3AtZ2UkwWk+09fnUFS/mBWzpbAmup5tVPPFYOpyPE/
vHD7DZU8nr938u/AP/llgBnSZdhu6lVoKJC8BTP1073cegHq3xwYtXg1EgNnznN+
PXhzxway4QVdijMJlw69VgDU5q7DY+qLUwIjmTNbDI5wYHvLZpr5cRN3sM0IU5gN
cRT2toajokUOP+09YvhIkaBTiO0G02y0OcRg4xAbEBESwI50otdIVylD9lSp3GkS
VfHGdRF49zFO+nZSC/oL0lLCQbZNAsXL0A+L1JsW3feRgHofMbdfiXCtZ0XRbdEV
+CKQRwFdV++FT/OSsvw4/8x+mbOfrdHXzyzVv1Sn7Wdrvp7LrVcx89X+vJAtClnQ
YKkVNCr9eH5CLTz3+vrAjdjoJWcKOKsehv1B23n97n6CfWNGKCD8qBicXTTrHmKB
SfYRBmWALt9jrtKStqiPCYnJGdaqsFjWPvY6n0Cbjosw4gK+Xrf6Xws4D5ltT+MC
lh9j8r6S3EFIUzvLxn3RIpxvwedCIwbnqSAqR3zd4ZLVDOjrVjQMvW5Ozt2ibWAe
gM4pI6bEGuLnj4gGnVu9HslprWJoAXahlZ60FZluYmAd5cz1/AA5XgrjifDExNYm
KzgltTEcCrpQPVqrC/NGqYmVGBAQMxLrBJuibs/B76YtdwJhqj485cFfMQRojDXo
jBEGpGifiNeTLtcVC3F/qU8JuA1LX5Qi+hYDsXhqD5UUsFyZpwMNOF/gxpgqqoCB
PKQHFPKZiTEylof3GI5BaA5yO+R4bBKvZDt6Cw1YTQhJ7CX71GhXgfaWoF/TvAmd
B61I4rFIO1rZF5b9cSNJCSfC8ln9Obt6XbbIomHYtm8P4bUuSwV2eYt4HSWG7FZW
hdIciuhGBMPFFBrMKnvXXhXcWu1hO/jGsjsGj7EpbDyclAV6V7zdu0SaQm5oGqC+
IY5pgivZ7bTKWNJVsC1p+F9NlSUXR/R6+jmGVp7CmCSLD9orDVxsLvc3o7BOXxWQ
78V7Ew/USux/n9e6VEYlHkS6F1k8bJ4C3OQMrphhTdpZjGU2+KzYSNLha+HDrl+3
OHbfoW2Mmsw6OfBfk9vmuIZpltQVKSPzvCYEB9T2U83KMZYZjvQgT8P3qXvVZ0/Z
+2/fcK9s1gOPS+96teHjfmGw7RB3ZVjAgy8y9SpWuN1qeuliAaGKt/hhJQONVtOu
fDeaywAjNCToCT9Ohe6SLHaa68+UEupDzGHJbUVXqqypdGeeFErxz/l2/gdxnp5q
Rz6mzXGAoX9Yb9t1tZLXW87EGradZ6cQg3UzbDiyNwsh4bCwaUMzFwSx0O5465Qf
1O3GTowsXU7DLutmHSv1gz3oLrxmu497P4/XWMyhxvwb1vUMfTQBhiLdpghPcS3e
RfoXd5Xn62Et3IiUNMO6iCzoOk5MpsQwfwz7w4PW1tV+tD5BGi4dv7bFY/oAdSOR
742oUWuN/ehRZhJ7Ou3KEZH6x+3d7jzzZY3vEKm0VrSNDIwawLcz5ZvBBc8wo0MT
l0SQX2ueVsMtJafyaU682OVNqVPW6jevBWUW8JmI9Vgi2sQ0NdQBAaNxyOwxygWu
cFQdfILI1nAyrkrfuGpBhc1084yz85PMa4DD6TEHk81ky4dMb8LAVDBd0S2+y2Ih
qxILmRiartJDx2ayaWyr9hKRaWu6fb9+Qgc1x1PCX4G4/uVA6GCdixOAenjslMiD
vHVYC+3MQbAUoYlVWyunqKVWz62pyBMnXM6GrgTDW+AANwUA0zoLdFUg40xFaJ1p
e8/F569mRfvTeY1lcjtigjAl39rEmV5z8BZksCTilDcPKVmx+VUsNSTRvHZEUBl5
CH5kfeEYRWDbua1/kt66sCZG0S3ES0L0jjc6GvChNrwBove8TVbyu6fIvPHoWmdI
UchFR6cbNakVByM2sIosH1wABH0gmYO4DOZCB/g03QUTtTP7m+iG0XIOu9yKbSwz
NQ696F3dX/hJJXd6B/VtNlixRfaBLcmYhbytwg5Ol8f0aps9pltLu7KEMu5vcuP+
LeSiND943igGUbmx4Q/sjCHj2ROEERbd/0Df7pZaL37yg72995yZNf/UP3MRn4zw
KAfG7oWS0TA7faKxCJdqD7OsNwXA55i1lOuvEeQsWnzlMI6OgNbqpsI+yScCH+pN
58kPfo7TbN+62GvSfNQ5YWTeaju/t9i0nsC8zJGByrGkFIPLdk3lfmW2FOSsjHyb
LR7MH6wUdy8D0hKbO5r8+hJmlu6pVGw/lwQ/Wu+S56BTAuBOowlbphIKmul/ij6p
/JdfcFjCkCO9H/iRMZL1pFUAPtFFsXn4iJYJXnwWEJN6T4lFR3w/F7batx39+l4B
zJ0/KK0n1dl1z8DIGz0TXg7sbVDK/z9+SzgeIBY3SRcewTtKi3fb4rs3w71d/ZbL
5SSQIqwBKwayRarF1byvbpfRLUn6po0DVcTNTARV0R0en9chpe1EMl3sOtQx9C76
SNuDL2dZTNbZoFyKWPo8/TBtVnrMcj+SPOvx4QHzVz1poL5J0iGOm1ZgqHU4N6zk
rqdK3rkqH3jzHgajTR4jUVI42XAAHb9uztKELbr1MJvcnAs0FIW+HL5lQFq1syq0
2ZlLqivPX0xQulj0jGBhaNxSkdgQ0uZdz5Ta8a8UD9bzCoqkviAadg9zTl+fJpoI
Z8aPIabBItbyyAXF/EQauqxxaQXpIzUyXSWorEWx/YT0ZpqZIvSK4VBLhjmViFGT
RcMdu9SbYphNc0DdiAJrT7arU01MZt06U+KGLeBKVNgiOqAsoPGNFMd4SQDATYPv
yVy3ZSLo0Tu79CEZ8LfKy561PO14OtQCTSKkM/+A5bYlhY4AE/A4qikgIKNmP2zJ
EH94dENR1qvGZA0buno+P5oRBZvSYruJIyF/626czj6LZC+UtRszXIVOXTHZ2QwE
AF7qeuuIeLCLDPx2bVM3OnP3WwRX+ji97Mn174mBCy3taImYKwfyjf0q8gAZO3Li
uyc2C2WJDypyaCkE2ZByxT0gZGY+cxuuBMFQm9hF6wY4JKT/Da4orlFOm8r43jN1
CmUcQNvtRyTUWZByHrt8vlstpS+pWW0fQ8iP8ZiXeMAHRx6LplfOJC1VBPxK7Tjy
FJO9++ZDKNNzTbdrVpROgBOxekltTw53kuxXWTRhIPPlk4HQ9Taxz6ikAnTTyFM0
2N5pnmLiU0HFemsPqrbu1lpxVZoUwa27MIKSGsJw9QdDRiNgLlY5T1LeVnWpAbvF
x2DYUeRH/Y9RqbR5xeNfLt0MlpiqlyudXApEiYkrEYKQNHQCsJuKAa9AkD+X4Rab
7ktfgnIL3r2qD28HLo848QVGJeldFGTcfKHwHrjS9jHrDG3OY8JALND4YJyCRAh3
qg4oDx5/EWLrOLzv21UkQWAgFlmYexI5AKEGhrD6gz4IJ0WX0rpPrMOAwg/fsTd7
yc5iXQ6kXsL2lNtw+Yq4M+0uTzCHMUB2Q96QnaLqrBi8cz4GbHnNDFRYiCJV4ilX
powL5WaG0uDnQtH8qd1Z2eUYrFwQCzg1VVzAxbaPD6ujvCS8M5IFZ/SOJxFUmb0l
Yh9jT9DjL8bCGbpJZBbfgT4YdwLQWr4k/V+nVbVYUWFm3rfYgQ+GEZF21V/7VdeU
Y9uEKNZmk5jgp4G/4h43b9+mN95jc4c1VbaLCBRJVeDiHg4+0KY3NY9d/OFccUfQ
r0HFs59Vtu1Htoyyb64uC0wQJMUbklm9yXbjKtfoJOtdro1OK9Y2j0f74Rb3B1wG
Q1U1xpM4pAESTSadAwreLJuWHNX42C+vpUNzRmza2rgMjPg/aGMptwLnzZx1XZWH
jLUeC+xjGyko2NGPccqypzMAPTRewcBbKscUs9SVXL/WMLDurOJkFn4QlpZsv9mT
YkUQMqaI3crYLt5MkZxb9t9UCVIyAs1ZlcsWjVfxxjIEZFIRYPIk5zXm5Y4ZzsxU
vsBZY+t3otAaIH2s4C/Oybz8LILw9MYXaH9VElR/1oige396/Uy7DldsXgLu60hg
X/RGPGA7oOwXtMf72eGLW/kI2hpy0Su5ZkaLtWrWGmCyh+Pt3HuRNkEdmEA1uUrZ
upwi5i2QSxHLzXnGWf+opAnydMUKVUaeLZk4x+Q7PrxvnJvCnKKBtOkTvP3Cy0nH
HT1CHbP9tmRBqF39yCZ/k48DI0AINzUdNsneC5vqWo73xEsPSHQ8GuJn1F54ryXi
R9Q41hrIvCEy9rWWvtTLXpG+FLpEl2LwRpIVlB+tKIiJwe1OtHJzCr6SulO3a6fL
3SDUR8DkEZw79UY9xHy4Ibx1SY0PBScaSB6z4qm9FpsV2xjV33CBc6bXM+wf++5Y
/0xv0vNhaf/F3htUnA6SkrmM8Rp+L0ZtjywdeVNSpyAnc1FIoj/YHEQVoJmbjrGI
iTx0weHygN689icpOATLHkuIprmNr727UcnnKCQVT8ftm2TyK9eQmfZt3lgII17S
EcgqhMoqHIYCmWA6ZcBBBfkNP/OlUbZL75AC2QHcKlPFJj9FTGkTXGoJ98ntFEXi
5xtJM7vvG9tYDn2VhkpCDlGn8sbf/e57weUmARGcFH8EeozdGgX3OtU/jB5+ReFf
ceVl2Ybp06BbZilLl14YPS5ZoedOoyJQweewrg1NyGB2BQ/3MWxGWmDz08Oi4t+q
oNM9k1HIdujQGap1ST2tu7adyQB/nOyH/N83IeUs3alLTKsISWldOyyNzM7HUaQh
Eecyq1mKeILt3jrmr0Dt9WVIcOdom10qdUnvtTTo7rBssTIG5LFHrpb013kcrgga
J+xoOMi9G/LalhNq5lOZQZNCoGTkSnrChEP+5OrA9o6+gF9Fr7qralVjmFG/jkum
8y85Lxq2e/9QH8+YKE4uXZTK5sd7iHnCDCfOJ3DWRFo1QrwVbK1aRrBURK5CHPqW
ClwxPmc0gS0AfY+59XjfPsfoqP+T919mIpkVkFYFiPZtMXZkSdc3OIFQdtblep1v
BfRhrHmTfHL/OY/R9yXoe6xl9vg9rwU0pU6e/s7msvJZh2mSdzQpwcNEXSGhzQE3
tUHnIUmPi0+/eM2A0KHiuUnCAncZV2azsdzExC4l5eJ638iHHgDejBIPgzMG4GgR
PKbPUdOaRxaMUEFvOXhVejaIJr+xuxV6pQFBT/OJycsNsIZQTTTZ1JUglvMbLkdz
iK3r2ZtGSbU7bylryiYgDQg4IOtTRx9raFg3jRZSXBOxMN1f0sPfy6cERutsDf8e
hHEL8nEaN2sxw/aStYgo38M+3CbLXPcjX/5kU93OtIUEgKvRQfAmd8uMx5uRq5jb
9UrniJM5xMMC4/3fd9pLyvt5VNV4fbUv5SRwASVQUkL99E6IUfstVZwSWDW2z0JL
xxbfH0uPdotFLTCueSZZTd5naTQT0gcVy5AprpiBvx320HmLP5mkkEXYfaHDXNuv
udJl9WieUXXO3zhPA0pOd1S4pPf4U9/JlfWnVU/OWJbU+tZ4QW87NSQNplnnOnAQ
F/ARNxGJEUV4JjloU4+lYuZyc51Ead2cB+vRaA5sxRNNT4wp3YFLoMDZg84chyDN
pSbVCZqCanqVeDQ+IeqFfxlimBF5vu5IYanmWjQeBha5wzyD5pNLz0MrWfCwTScV
cyiq5Y6LfwKEpwp7HbIKvCbLu7ENmOic6SFO7NY8hYSR9szjrtpK9X8tc9XXBJqh
piCn2Jv7tXNInZc8Wr3d1+JowPJsWrL9NqokOXztdUxZsmjM+ExJwCWuoVVZmnAX
OUuT1PC5r3jJO87zctMIHM7U/0OPYsNWtQ6pt0TL5quUmuxhrwRK0RvbLnJb+x5W
0PNqPSPAv0pmRxC0KYz74ssvnlsCYKTRyRjFcglEoqDr+ryPoHwRKwzCdRcPcV4q
c/ASYoCs2s7isXF8xX3syjVbk1xdAaspENstadgmBJRzXIi7+TbCiuxS/RwivnSt
zNbro+TwT2dss31bvNTuM7BZLMWzvQt0n/pUbeLEjZO8G8U0sDbGSLLNIotXswtF
bbrwUKDMy+rvhn54d1DjCLKa4kg7EYDu+EU3jdS6Nzm9qD7JDSe5yEx/OS/M/s4r
6vUqO5E2wQ50zVLzSg7HtpZEn2ns7iCgYtttY8+NnKxRlM1dHT3B//wzLGC5hdA5
NcfXH+Uh30i+APboDKipmR3+IBthP7rq5WMlj0EEiCzy/bRcQXUjLS1rxpoHYDG4
R/4nyTUPim+G3SLFT+RBwnb+r4SL+a90CQJFMn0ZaE/xmv+GM4+6wj3Um7xmUpGB
6XQM5i1PCdJs84SEcejiU9e0ZIaFPmUMajC9xsdHvZZqCuHYg1nz8TjJbCpJz47q
EhwRfQXGqL/p5eUtieuKd+U676JeyMV4sOfVey1QlWNZ+KhRAIPbOGFZ99pDGyKr
74QFueFZvjh5xZgpEzsemhkZ43WxtV/svvIE1M5eycQycaRoXECX3ANpD3zeeshR
pNIniufmyVgqBW/Vt0F5pEJF9/fUT0AI2TjVif8Kt6StQRfEEjSEezxNRwNEVzGk
bie5e0db2Ni/3+v99tVOvHa8+zBYRDts8oNo6NftdpGdDANIZzbUWI0zYBvA60Yu
bzLrg/NHkQiucNZlw5Yd3Md/z3t/s8NFs+nu/OtCYF3+PxqExEMPf+OQ95tFj8hp
UqmDQRFtihxDeKbCgZrcg43Q16qh9sTVqKsvgsIU2Jsh3YMM4viDcWQdyEYD/Aa0
SuHRXD/ucJDiJ1h+D7pXOzAOC13NfmDl4opjQt4wwJwIS82VqzD8WNLlfyKjtGcg
raDQgkKH4XROVY2Xzd7JcjQOc1BnkB7eBhh66obD2LNk95d+Os4tPOaG5JwRXlR1
d3YgAEzQI+Shc1KyNb/3Ngwro+FCMSyxm8yTwex0QpE0vQ9f0fg4VEE3uoODOBEU
CK6ciYRh20dGjp7DZN+bsx3gdUvviuJVRa5Mq2eJhyoEyca4UGw6dpZaHaO8ptab
Dwp0QzuH3+uKAbXPlTqHJOhaAgBkJjdUSw/fp0RcOE7CZkgjF4lJmKRMfSNOnbAJ
mDGrCnAn38FZIJ2oTE0/xchJ1E+FGNLQoeEUQ5NJmF7LWLyyE8xyjpYkRCW8DMXo
WTQprr0pfngFMExDhJbkDmW49RJJTdL5iwTNQOAO/maaJR/Reu4Q36+1WuBb21v1
C9sIsFVDUvadlfXbUJVpp3xnvfA71SsIP2rAKqEAgl8lnLI4lOLbqQr8EGQZs/GX
bX/w2giyNZUJuZUX1eFH4LiIWGBlNkzC4YCIEB5Yb+e+iNV7Ywz4r6yOAoLOvHBs
RC5a8N6mntnkTUHX6jaDO2Vguwfm1rtdVsWODKahL1WrQiSmzm0RwpIvsU60+x8u
0Q0f+yaLwE0OF0A7M4Q0j9yrMJIT7WPMYdi3g9rSlA8E4bNPZeg3P7qM/Fqx2cec
lUoskn2YTXYLzpbIuCQ96mU9VkHJYt9kSKraL84cBTnm9eEHvW9JdzooQLv1ZN+9
GBMFOBlXAcbAdeIm17AZQfrY6MsbKaBvAXEFTkmCo/zvdYFtcVxJRBWF9QrwZrHn
eLlcxsp6iTBXfCUoRZfXkwAv8qIvqNzJ3LVyyW3V9+e9fWVOhiyN3B/rrdxXCDAd
m6lsyZjEMm83rn2dciBV0fqEMralWAAQ6kjSdfYeC4lAlEAWAOQqyelVCUNWa0Cy
RFxkdsXIDVySA7Okabo8lMgeT8ZaX/KjuSOKR9kpgvVU+DUhVoSsB+FxZZKOKvrU
+qVP3c4bzS/qvMN2xuVualr40T5me77+HhvIABFfzCHs/7kVfq6VplmGs0eSOAAx
Y8jVGrnm6zB7oX736pOML2xh4tFR9dWTQjans0Q6jWMwLH0BtO4k0JohAJbQRNAw
H2OdpE3DGhUSFvIakFAl7gjWUq2xMZf2f+qZKp3IoHXtNqm2GlshUHEPi1zF/Rht
R3X0bC3nONlbpIrYKb8uH5f7czD2JKVNBfupV5RCGtvuJSGP3j2uwSqEhAtOe38Q
juJVWnxV0pQwV0EfUERBxlu1wbgDqkR6OzpE2rB4u2pNqbkB/zgkt5CJQorHXOPp
xcRQzug3v9Y/cjB39ftkqD8knPRhva0iZTrAHAXgcBxJi2qUfEmS/mikRMDPNcoO
5caG6EgZ45MGw51pz4TyhPjDinMqPefAzem0ldJkVci/kMbps08hqTyTNgvj4cXe
g+cZQedf7Y6oiHtRcJ4FHVYfEwoQp/Nn6KDKO+jw3e48KKhcVuTp13zeb9KYKOuF
BNZfTVm1Y+DxSj5pN4PQKrYcMlHaFvXysD4R0xnJLfLjspMt/PoSPNFXMzvJJEje
f8vOP3Bl2qY26KSXwJwS0ucBPeL8o8c5/M6C2cc4uxbyRM3FFpiYOsu55Dmxjgiu
nsYxLw/Yfuwn7ppvekobwiVxjJoLFxSbUOvI9o6WGn/hJqwBUsbE9UXCru5eERZ+
3CFZyhdhqw9QE3x/F3+C01RbbxUxDskyN79rKY1FO/rDjbznF2cnPj2QAz3i0Xgo
La0NUED1AO35XwPpzJrqaT7kkdS9AzCdRR3kVOOzXRva00HuVyGya2ndb6qg7Br2
WlqavaHSZdYyjr6M/zlZqhNWSZdC9VrE4/DbeViGzc9q79s+YsXmPGYJcA8FuCmG
MSsddRleEwwktfdfkI66IZTFE3/BVcDXA4u7AMG6JD4xnkyDx3ki5ixEw4Nwb0Sx
Vgktet3whtn0X0CyOiholVARuMTVcECUBrCPgN4Ls+B5ZZmzZz3cj2XmZpJ7pwdO
aZyzsW25TajyC2dHEK2Xnk8uiW1RjvRUk45hTsHbzKlgSYpSfcoQ/NZD4NHtMyFH
7nKypjdANp43nOk0DGRYnc86Yoqd6Yll81GEG6Ka4u2nxCYYZUaaMRq4cqN3eVPZ
Oz8DqzjB0MAPP7FIHHXzz4r6Q/jjjDuvOvEwBWpKqFUZdJLkXO7J+K9XmMU6ZpKx
obS+aykvTvIznt6Ks7s6OqR06c5Y5RYNd3Gz2x36b0uT/ohslEO3mT3M7BdyPJrI
xZ1D9JJRN40M7ik3gG++Q97IyeB209iVDGQBZEDBV/zstf7lGYiv9CyitqGfYeRg
+nbuoNPumA8p/naXxroGlh5Ib7wt99NMrI24rPPwORbH6TyJU+oydoWFPAc/r4jI
DUVcaQXCr+h7LTBqGoAnW9Z2G8mbrjIUPbAF2aZ109WTkuskiQi3PwHwZ0nvvY6M
AeeHRwG5tGFML9+4H1hMnLpmL3AINm+/5n8RT/ROXV7bJQrYLr/1UOkqrnl5kbo5
CUCl9V267o34Jm+caumKcAuQ3PNtyc/e20i10YGm1IY+iCXo0s3pOwR1cxnDu5rK
+uHyUOsPdoglzMy87cuMlekajrkQ0JeLqwEUqyPlMQOfrW0pUhkQDEp0jMuD5Zjp
Nj/VxgU+7bVuE4lh9sv+5TrjhrsL4UMcqBZbzDDG4nfN8ICdMdyX19KNUXTEZTDa
eT0wST6Dw8yqAO+yqjwQoNmszg7CCn7qTbiiU1sm5tqvc+H5x897ExqWspskHBrI
299LTNDpkJhiG9uDkCDXdXTmGXI2ljoeCTE8aXLTqVRlfMXGfc0wzuhlLIgyJdw2
vdZp/XUXmfN3/lnD+LXGc3qEsXjeGpU+Tht335qhY/F+0iYqnY7FfdDTLEW98l/C
rX1I+S+QtOKp05mtG1KY9a2rywrjW7ahrzbJdb77U3iuqDNtktM+bXVGoL+qrlD+
5PPKUJOlEFgeS/KplsP0GmvBkUCqcp1FuSGlnDvWVkuphVmttrCMrooGEq1FC+zj
gUZvovpaw3kzfDmWU0bCM5iJaBc2EpafUhyIycFhXvOvzcFwf/3U+c+eMuWbd7hI
97K+ytSgjyZjMpVcty4fO067QEEGC+pSlqdVIG9qh6WKEKBcE1PrQo16cLavyK8v
Y6zj4cPmvAHb7eZYHrtk+b66qjdKwt9qjlVU8Y2WJfW3Axh5ZUERZWkjdYRYZLd6
Xkdv6arAjvLjLJb+eInkkXepoQjhVmj5ugcUaoFmr8ZW5vDEwSTUddDEbFOKmHuo
PdwuZ46+UznNc6OyUpDoJqZoFVh5JtGS5C2jGashNS0wU++PwEcorLToLsVay37Z
5ubUePASFlosyTFMtzeEcfA5rfQDy8KEHO1zfFYkXrhGJ1UbtnTbJ6Z7nejzp7dd
1haBMwhgjXn4EqmFvXAJSdljG7NzSxVPmdWhr02H5hZr4kKCjT80aVIukCp1Kzek
G/kB8QRwwsJAF1S+2TjfXme4VmZOyGdAqD9vZuPQD0ctl8eI7GvlejDUScP0AR/r
SN5AW0jnOiaeJkcTEFouI7vJNlrWcHTxHalXFlljXnJRMKvUWochpQu0RT1yHh/6
2Vg7mzNJzoi7RWG5QkDiVXxFPDWVB/oBNlN0QrDelOEYlVGSXfTaqLinO0GzEoTn
75bRcnUj1+SWtRrXVmEGLaeHta1YCdTpmlJ0wAtkkEbDZ9VyxUrsrSydaaukIyXv
vsn++eNBqER92wEdfKRNHJb4GBCFiclccwu8pNexN3V/E80sJOBapWjo3iNuWc69
KdBfSoFnwMKJ05VQ8wUsjGPO1cEzTBpgmeYrbTForsv8leymGYO6nRSAu+LudcfN
HD+LCx9brO8UoMCeP3V3sfJDxhAhr3jIQCH5o0QEu+TJUkbF+TVIKIGs0/hz1g+c
0JH1GxDYUNM2SHWlx+ea9UOWaEvES+Vsk1E50rshePl2bL2+dZAqZjG2TNReSKez
E1cpS2N2NVHHEzZ300cZx/xQLlC3h3ISXWpLWeFf+wQzbiQ4eWqDfUqkHGHKo/cv
NW4J6E74NmVBqG6Eto40FHkuvy9rrId1dKThaVdSsXXSTEu6HIpwDdN96jyfefqa
o+j57p/g6g6H/tXJB+ZYtfmTUlMm1RORXdYBlIHsrxKCoU58IkETWEstMV+1Wyh4
Dpk4ygO0cr/YcSjvP7dxySTbU1Qz0rwDxXb8sqzz5h+9Bvu3Z0fK9yyt41UuQp9v
BATx5EH3nSFYMMeVvQgaX+PFhC6PcE8UvKNRx+D8HkyfgdkvKRt6HvU45/cm43vH
A20eXfxEXF0oxSy9eU6lhIepSE8DHF6Gz7RUatVPsWlbb6NkI/jlk1/jarZb+f8C
+WTWg7A5Ngi1BY0kTzhwkdIKiPImBucDY75U7hKYi5cfskt5vDw4GQpT/EfkeDqy
NNS0yQs1DTTDOaDrpe7rJHlN/insLybSNLUfGyRjGLdGtwvrgXnyadDpSY46H2BA
6dME7rmoLFTB5Cho4HaamKeCpeCAHg6pnvZ3/pEHuMdc2DdvCZ8XAl4nFsqjw3M0
1mTFzmbEVftp17JHJbTjiozYO307sjhSKUpOrDlfMSx3LXlBGJ2PE/fjD3ZOvUGB
swjUqUppqJMljFkejuiaulBuWkJJSlMGxu4VQBw5c92TvTWL+B0dYs7W2FLifbdy
0t85Lw8KWXgxbTKi0EVpVZ0DeApuvHfGaCRCS44YilBWycWXPkSQR92i8S/0rgGr
EB1bAoBpBuU6w/lFtW7919yMWdoNKmN1a5e03Zu2xLGTFvw81firAIylQDe7gOAN
SMNjGLUW8CM2HXzxoR+olbHPN5/VXKCpt5VTKvMoFljL6eWFjhCCRxcNMoypkTQe
0zuohT2naTZvq4jKkFDXxwzg3ac7TJd4PLvxww2Lvgnt738SNGuBvxpQIQwN4iKY
KTPM4p02Wjb9Ehgvlq5Ag7K7zbSiQFRfvtM2wCHrLw4AO3FkZvGcVzpTptL3/ABG
yOoej+uymnspt62yTyTXg/RvB0bpphn5+uOh10nEKeFXODpa1Kdufo61mlGmaFjC
6ajWX2JJJS+RP03hdgJZAeOYvcXRFEn2vX23MwWAb33gvsIpS7SLrRRX1VqcPIHk
2Cqbar2gRfmBcZ7RRnvdpZYBZANO9r2AJsJyQDlT94Z1nejLw8/7V2LKwuKoZCrt
2vC3S51GrtH45qeyw5jJXSu5DZkJRHwsWIwIRHjGd42UjG4GARL/2kXlTzULsjKO
kWYz3YZ6B8hfdrDxWUZazk7pznuWKgEmtesnDESFdwQiQHfnMzrmdCiOqB9o5v4U
82/TYGX6q+Xs0Hhb7MtCR1tDMz4OsDEzhUMyRjZJplwC891myBTZPYV31xaucMZY
DkmPBx5MAQ1kyGEugnkeRWwFbRU8BHv2EhbZLdM6OyT6PbuFrG5HC2xV5w1YMjM1
0A1/Lt7mT1aO6JV3EZyf1Kg/2FhgbErfIDY5/+xXV3P0bv9SFWHyggKYT+O+pfdr
11Rgm+P82HuP4tZx/pZ2AwzgB1OFUF/urFwTe88+JnuHN/2ahfhD3mFzJdq7dCiJ
SMLn/49IlVTXeV5C74tkEZlx8odYsnJ+MRgc3B2ImDvmn9HGyz8hGnfRxShCZkgS
gGWE2LFRxqVL72ggjSSPQhFvrJ53HHm7hZeeCsTC3LZpssbKWFiuEq3wH+3hy8vq
3H6XWU/zWWN1xCsHZAWtqdU/sv/YHwtfUPEO1PxDe7zMOo9/CYjtI8xb9+tSNmK+
Uu0aBooDcgVkMxf0OSxLetESQXnqLKZJkuPoT2lHxn5ecmFL+n6HRtt1LWbX4UC6
u5LnzIPEU+hRMplqS7KUt934IozLIN0y9jjoX091V3E1oppq33wV2mPV5LHqItIa
gHU4U9dCaJelGIoo66+jWdqJyX/5092ChFiMxf80VNyYM2VLIna9Cp7Xjil15p8L
VG6zC6/592GOCZQCKy3YK94VcKE9UsvTij18aJ4+6Mc/4rD+J/GAGWnGdsSG48p1
QgcuWwLcYqlAQ/P98rK1zt/cDkjV0mCM04jKsqyGvv5u4xx1MBpYwDiU67gkZJQa
6HKM7jZdNo0h4U6zrbyMYSuSW54Tfm7mYdezWyEcmRvnFmA45LTl1mxEQcJwiVXm
XAy1zsqjyqwJzl5OpiKqVQo9awI5VGKRn7pR5QBOlSMgntEUT18yKEdHqLKpx92H
bt4ekOSb0CmYqJPGV++KAx5ZVs/d3aZ/1qWmZNCJQiJiygLaqyFvuZfSNyUWLJ9U
YDZj3GGthapg4PbxnkyPxNmPf2zGzmUCng9eAlbNbV3bKckmsTtkQmOvt62Dz9yC
D4h0E6Nnc4omx/8fmN45GgklSigcQmxv049MO2AvuV2ZDlN+XGDvB21cgFoNHQ9w
ZQTT5fQCUpWG4CRKzfJE1TYK9gBNUZbMVFB5BEgO6555oav2NC2hR1o4MeztEtqJ
HT4OQ66l/HmYWVjWEvXBhnIyXyMZqDYnT6FYvXsRCnhY6GLxyCZgUqDdB8lAGGnK
plvTbgzWQPUHve1+ZHAzA09I7YjcVCp7rfEc2FTpF2oMpDZp5ATC0hLqJxjkFUyb
2lyjqeMO1wm8Is2pb4kIddVEBcj1jBja+mOuxc0s9krheCB9iE3YvZEK9bIy33Gf
NL6ksGVrFFkDRiUi0B+99oXDtpxB/dkK6+vCMbIbaq66U/GAmC9i/cOBxlkdmGeG
ZPBR8LsbOqwpH9z135toka2b3pHSplU+biyD8x5Md28vcpIvdwPc1BX6jEejfa04
wh6q6rr2qFO0ObhUfa31ZHo9HnwDFnfCSyxxCDDzg40A6n3rpkQhN8+6GAaNfpbU
5S4C0t6MX2Q3Tc9d1VgW227SiJOVbnRRh+Sntq/ngPEgUqxb7YJcJVWP8esq6cB7
lPbcbJlb75i3OxdXB81VQMGhQVy34Q8VkQjFVmmMSNgHgf9agF4OH37iC815pCOQ
WmaJ/9fQDFXNQTz3+KCzkrnqor6/W8RGISLt+p3C2NXI297fgcnzZS3td64bCTbT
4mCA8RbofcX5PP4Sof0hQboGf6mpsR33U2fMIiCosFuLrw8ua43VaaVe09JdBOxx
Eb1D7apAIFneDUJ+FEM1e8/ePvS3+kF0gixpFev8rFYXhdInP7m+A+hzgeW30T/0
xgZL1TnGsPSyW3TG2lDpxg9/que9VkK42aJsEpEp4FWEYq5TiA7u5YVNcUrCM0Px
ZuiygqIDG50AYLfdMUQSAHUlFxh5abvosSsFEGhSBb2rPRg/pg9fNk2RCMkBj5nR
jTjSs/YEUZ/h1L62ri1XIDFNNYhl0lpuELQV2Hl7Ui1bqJejRo+fMvB+Qv1RjEsY
knkKwzcsiMsTT2Nx57bqDvfHZinwuGAjsLcaSOB21RC8GEAq7jxRm3zI0qulN042
i/t0zX4hYMiAkQl0GBcTcEI0nWpHtdTtjLM46bVfXmOvLyqikVtH5w/d2je4nSpK
qbIROugf9IZbfIg2jOhqT5XltqItwtuzRKs9D5o+oBZFpVFt6SDkhUYvz4ZQk51N
Qah10HiiY25eYSxCWWSnR16in+GMRM6ekCfUyaGeeOiprzPYsh3SxaZyXmc1qTzo
YJfq99FJHdPcHoozKCCUjWgT9HQgt1qPijdOtkT1p11LRiccbvujDqHml1ZYmdcn
LFg5n5VvRM1l8B55y/3sehSzyFQWhWExn1VfyDxPbuyjBF+S6EdJeohTxJYDw/Lb
aYDdRIeQZFIxBB+oV7zCExhp+iyZ+O/RbEAy/nZ/+0gEl83NvrUYhYFAPyvCZ5/D
Y785AyinHX1jhLWxkf4sHHqUyhMg4hQTEXhF6d/s42gB7ZnAFSXf9v1LdzqUCrw7
nY5ly61f7qutDclZfQDXCOR/cuWzAvNwbuTdYZs8DNbOpjuLW+8JTy263aputaFQ
KGEiwljdY+F8xrGbn9yAr2Z6+eZfuJADKxZ7q1NbjPAnHT7HgObue6z3/c6Jdodt
SueJHHZw4Ilc9vs4T1NkSQOWJ3An3BQ5Z6o4BPF3KSXBj4IOTjyMrs3Tg1+ruota
yt626AtrtmX+xT+Z9xXfMHtYM7xh6s9HIdMWrrmVT8gzsCDcv4QkQLsAEJ5Z7nVV
hjw6CB3AvkR/+nNTze56M+pOX+I93TrN/2v0MgM/H3/D/brH6WBP8xvIXcB8eoNh
A5iW+ywjkj6CIiHTA0ldAyfjD7waAFunPJfrtorl8wd5j43ad9+F0igzZAbQnVXA
JbWBuXQZ0Lqx3Kjc66USKwdQEWWgPp2K0MNevJOzUIzw/XfgOHWmUW4WgiFTOaRP
xU11wL/WuOwqm/69MzO4Ww==
`pragma protect end_protected
