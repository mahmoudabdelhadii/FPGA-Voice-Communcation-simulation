��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��,�y�}�ǰ�=4d�H���`I"��W�`r���T:tB�T4D�m�)�	1��I�t��
��8(�8t>s)ו�."[�漆���]�~�]��;�O(1#5�-� 偙O��QZ��~rL'�x[�i,mׇp���O�I43��4d�,�H�����SN��d���3���r��m���̨T�I;uj2Y� Er�*p�Q$Gm���p�V�`�2^���,hz�<p��l�Bxt�5��s��\yq���#�@W���f:m��T�	,*�񞭋����_��㧋l�	�\�:��uGd��PǷ��N�I��_����Tuv� ���us�(H�~�{2H�:Zor�Q	#%�3ˠ!��iS��95�,?�.���/�F�i{#���Tp5����Ҥ0{%���2vpn���X�����@l����3dc�ק�3	�Ed&3�ZN O���z��s�yxӡt��v*}ԫy nj#��lc��m戭k[��5)�A#�����8�!�]�Z�s�M���t��w�!��'ÒE�rv��Ϝ�c@<U��\tq+��&|�&X1)C�����r�A~��B�&�����s�:n{p��͠R�X⺂L^��R����c���f��J^?��ܣR�O 1�rV���:��T�4���AD����˩�F�w��)Dm�O�b,�a���1$��c��7t[i2>�ޔ0,S���󧇳Ϟ�ᒨ�-��}�!6��Jyv�醊�^_�(�H�(y^����o#����X��3-�k\8�M�T�"`R�DF6ȕ� �,5�;Ҭ C�k���1\������k�t־9�}���� ���QHF��"��t�9 ?��{E_�7��!����](�S��0�q��w�9��=�i]�1�GʦȪc�W�XC�|�$��}q�6����zf(����լml�dz������*�eLD�*�,�m�]ہ6����D�Gw� �g��' A��)�m���b��ӎ���o�6ūvO��=�W�������}��	����z
��z�&�P�K#�^Qץ�_������&�)�ٺ�u#uD�	' �/|�qf�M&P)�tL�x�?�u�����ҽ�����*c"q/�\��YDl2n֢�vtX��Q������ǰ�6K�gVL��ο��Q�������-�˚e��"gb�_� L01�D��ثU�8-��Nw�@�$[�>V,���6�����=����{>G6��v�����φ+Y��	�d�A��b<�)��Gp���k�(�vWu����!5fQ�s�}ɘ���ۇ������4�~�y ��;�y*�]�}Ox$5Ǝ��)bNA�%�o������;jE�����dU;J�5�?te�;fƵ�L�诺w ��˘Ko��W�T�HV�w��s��<s1�a��^�`��I�PM3��1M�=(�1�Lg`�P·A�Q{�T.�9I���p70��:5�c噒�.���r	U��բ��2��I09s�m�/ah~b&~S����}�0L�Ej߿�ޟ�j�����k4B�y�g/:!A'����)z6��.��[N�ߞ�,!`<��-�'*�ȑ?�H	]N�,ꥀN��Č\L'v�m�It	�%/����r9Sw�<lM�
��S� ���l_��>��G��!J���D���o��'�R̾)]�=����}Ȩ�5�?��-��߳|P���{+�[l����m�_6�9�)�Џ��x�n�M���Ka&����������!n�w�۔�4��~"d8��ad;O,4g��x��1����ǕI�{f�v>.����V��h����=@�+ҽ�|���Ox�*�2�o��������q�C���{ŉ�� ���M��	�c6Zs�GW!޸�o���zo�y��_�U�A��sL�jJ���ʀ�bP�����y/}NMabU�X��z�J�C��z_ΐG"Ec;ŝ��R������:�j�;W�[����Eb
��X@��y�T��L	�&Gg�N�$U����:��L0����*�E��e1
�V���65
��.lL��R�`�x<o7�����N;p��}b�s�����	\��Pz<�W�-���灬����g.uu,.N�UR�>���p��g!�TX�RA�z���q�Y��|`%��Ţ���4:�����7�3�7��tr��Id���u�}%�0\݌%?_�����A�v�2`�sW���;�?։ �M�H�)�p�4ܾ�?��/&���PE������M��-K���T~zS=���f9>�I^֐�]��d+����Y�����(�J����ڑgnh�5:�k�������H��e�xP=Osԝ�l� 5����e��H�Y�HG#���1�7Ӄ���[�<��J�P+p�2�] d��@X���
ñw�57"wR='�е
G�4��K�;�n�ăCr��7�^�R�H3.�MR��Q����(0�g�^=��bb�:����l��=�/���D�#���0i���tR�|�yh���5M�nt�"�>>Y�Y���a��%!�&w�7��5 \�>(o��`a�2��w4�M	�����T?u��Q�	0��{�*�f!� Se�˲OWq~ς��G�亂�Ӫ�����t��$Ԥ�f���E�C	�A�3k����A������.΋�q(�]<�?�۸�h�L#�+T��I�(��`�M&����,�n*l�Y�ka�"�῍`��y`à�i�TјԺ�'�JA�g��i1x�U��s6_m�T�+����5���R��[d�\�]���,ju&�I
w�u��j�r!��߯k%�9�6��	56��+�<�m�,tP�;��鲉�t*c?=��;�a_�Z!7��s�L^*EGsx6�=�2ՈE
̆�.Gw�CK<-έ����`��hNi��
a����j M��F�i���xP��B�0�0���u��ڢm��LI_��!^�Շ;b�
�L��۔C�,��`�����/�lW��m�P�-�t�.�2����`��qJ��'�
��H��F�s�}��`�"vbkg6�m��e��"�E+�Vj���t���az}�%�I[YZ�[Ez�I��)/'̨�T�ZX5�-AY{4K��ҕ���55�J��¯��;�w��� �4��������MTރ;�AN�J.;FΝ-C|D�f�����w^�XuTM�7h�=�����u�=J��'/ �y8Q��R�G�量i����$��lKO�r:ӕ��}9^�� �[��2k����V���< 5a;��ƳRc~�5tg�R^����Vs�@�cX0��⸒��%y�p��$�Ԅ{���B_&X/��oѹ�3��(B�鄪a,�$���=}������e�G`��w#�&�²�VGv�qthܽ|S�)��{5J;�3A�tL��@����JD#<���9U3�Ey� ;�fJ6��l�K�x��%�����vG:$-Є�h�91�$jGi��K�n3�ħ����L	B>��&Y��S#����Іaa�=�]���˞p�1��z�K�cdpE���)�hQ�* o��j=�i�y2��g���CH�+0�@5�N�4	$�Ǜ�$�|�'m�v7\U�W��-?�SOӃU��3 �8�u"���{��m�g/�$���c�s�8Ή��(�8��t娂��F�}�kI���-h6;%P�oI-a���6���}ϕ7���ڡ���������n���Sì�4!1��`
�_����jBgmj�~�v�:CyeYu��a�?���%:�,9�������N��Mߪ��!�����x��	�>��Ä�n��.�h����@�u�-?�?�K﹤�I{��T�>��y	��UX��۫�_�r�+��U#�x>�\AC��v��.E�N���c�}��.�$&�yd��q���B�ժeg��4�vַ۾�oN�A����&�%�ܝ*H�֙K��3 ��q�jpo��տ<Oz����9�ܝ�\��'CC[�֙��e�x��'7���F$/�Y7�b�h%1�$�E��6:�w"�A�B k&�7�x���m3c@}��m�X4n&��/j�(�d��f�����HP|]hTႂ3�$�A���v�E�%Ӭ��GĤwG��;�Az2~i�c0@���U�$T��$�\�	f���.�J�)\l���_�ؕ������n����|�����)�»�p���PQA*��/��o�X-�S���[��	U����8ŵ��5h�<���#�$��,�3���k3΋t����Q�t��ϒ�t���=��<a��� �!��,�t�!NR"$#`�H`�^�P#,Ȟ�xK0�z�ҿ�.a����G����~���7M�3�RW��;,ɷ
%�DA���:��3C�l�j�5������1P+!*���Fu�*3��sa��T��M�~�K��oY���xoI�!�����Mk�<�;F�6=����*t]��i�^R@�#���������}��XO��s(�ׂ���<�X��U*lk���K=����W��8��
�W*
�|z�H0&Ef���2l���H:�tmQh�
%�A�����������ka���=��?�y�t�\��h��n)��Ԡ��	2?iO�r�2kӭԇ<��d��n- ��S��%��9����+�;��!&ٺ��~+u?�F�	���J����G��A�Y���d�3I�<���C���~�(o���E�]'�9��P$��'s501� \�@�P^��!���kD��Yw�C`avU/픓�$(aJ��Pf� �T�y��pp�]%�c� P�(��095��}�Pp�W����K0�$��ޥ"6𔞸��`�T����MV,����,���'���/��)�e#v�����9�Xjs��p���m])�KL��x�A������ڇ�t_ᶫ&�Z�$�r8�_��P��=G�2x�2b���v���]�ZR�x3W4e����6�h���J���Q#B���ȿQ�͙��3x

܍b�eFp��O�w�`�8�c�p�Q.dD(�X�6=����b�΄��p�dՁ��>�E<�#z�'Ԯl��cF�v	�=��\��&��V�}�C��#����4�B�����߮?L$����kLO=Լ^���+X󤪃d}���&�v��zn*נ�
/c �U�la=-�:Un����\���� /O��� �� O�Q4��*� wr��4[XW�5�/�C��4Q��W�&o.�� /+pYT?��,��r�����bl���H]���R_H!�Қ���.��F�l�E9��&������>��Hax����(�i>�N�Ro7Z1��$b\�!�%�-8MQ?�6{BҢ���DKW!sw���̎������^�ü�'5�t4s���r��9�l��k�=����4jCؖ���RCS��8���]�`��櫿���Rڥ�oM�F�U���3����pB
��6����Ϭ������@4�+D���nO+��^�rG.޷��l��[۾���{�(9��x:����(b��4-	L3�~�zi��-�+�|M2�h�_
�b��!�)1��h�tb�P�\���Gm�4*��H�ܧ�/�~�ź�m��3�Z	���� 3�杨�a	� ��X�ep�1�KE<2�&��[Ƴ,�!"Umh.����0#�����j{�z;P)K�-TڜM�%D<:<���R|�D�Mr�ܨ�L�pL����z���g@!���&LM�=���|`.�#+ʀLR{}"���I�����r��s���ᭁx�j��P	q8@!I0�3Q?y2�Q
�2��X<��t���ŷ��d��R��C.�Ƒ���t�3t��.l�1���c������K�/J�#'I%6 ��"$1� �L��%���!u�W��C��PQ'ۋ �H���(b�#SO纤n����C�q�r�������J��
�92H�nTGx�\��G58)0 ���j����2:e��XǬc��u˅M8�X�6��n1fI]�O����g��Ɖ�`QPx��	��P��~ ���Ý-,�ҤF;�4���I��l�"+��k���S�V�A�"I鰌���	�_�I������Ơb6��)�ڸ7V��]�0��\֒�ٛ:'�����jF'�&Tu�y�o�[���x��*7���թªU��<�i�� ��u�q���\$���98ƒJ^-Y�x�ׂ2 m�? Xm1��d☟J<׶�i'�f�|�v�~��I�����&1�F֝�d�v�R���`,b�}��3��	��׸�vƵ0�����z<-.HG ��GYd��C���$�|iZ�쩭�i��'�{'�)m/[.6Bc	+4�`#��f?�h�(Lw��I_ �b�!�>>���~��3��>�p[eS(?��!��j�Kέ&�dj7�T���\��ᘖa����#�^�/����Ux�W�����I�s�Mw$�3e9�?z��z�|�2p�Heן����ZANV$�p��X���y\����Ŀ�ܾ��a�S�,\���R.��;f�f��,֜z���҃�Re�#���3x�Ι�A��z�|4fP�#��k�ړ���MC����1�5+�&��r��a�
����ll�MO�F��;Hm/V6�5����̍���Q���?���Xy�o�ɵ�����&���B�^;GF
7������?y��YԢ� H�,<���&���A1k8�r�u��e��Q����CB6Cz�3�7[dmD�H7��c����#�V��}g5�����$��c�?k�P5�¿��~�^�>�A��Yd��8��3�S|�` z3�F9&Q���ƀ{������~�5l�l��Yo���+>����l��lt�\��oC r�z��<���׏G��j��\d��Ѐ�U� @������!�n�[L0Ǚ�]C7�P�Q@6�����twŎ��&ҝ��Пr�+(%��y��7f\�Ԙ� �i��)�
�H=Tu��$�ڹ] ���P�+����Ae�|*Q��y��ꁏkP��J����y�e�]ʂY6Z����/��.��2#.�O۠fr8Q�(h@a;�R���J�4p��<���:x���qG��z�����u����z�w�a�5@���G�tSj5��8���J��t����]�(=�3��5�-��2���f#�~��χ5`|����՛���	au3<��ꖜ�pw�0�V��;�9_\w�����^Z>ֺ�Y��\(�j�8rHc�=)���R��X7M)cK~�c�Bs?,���X�_h�iS%Rn&��<�"r/~-��h�JF �_KG�U��|ֽͤjA'S��5s�l;���>�Ћ��݊��8q����{��̓v�")	�*�i$cg�]���$h�EcAb�XÜo��O٘�A��4 �<��P*'���0WxmFjѐ�&��\[��sQ fA6(�U��.��׽�+�O�y���N�x��}I�9&#����,/�jN����V@��4_̓_0�`/"�	�k��e�r���q�l�X�n.}���A�	�{'���6�O�����Vz�F��E�,�����CH���f�c0���r�C~��e���?��t�W�\n�� 5�@&p~r���gt���������ɴ��*��3Vn:�˫f�LB"��Èh�Py �W��Q�9^֑7�$p�Z?�oދ��On�"��:ԎcT;�]��B��i4W�}K�.���39�hPħaꮞ������D�g���|^���s�z�\�q�x ��׏�s��=�'ym!�w�;rO��S����!�*���@���]��@��Oj�3c���Y6��ܝ�d%$Xh���J���9�RQ@��ky4�=*�a�6���s�'��U�|�.#����+3 ��V4M�,o��s;��}�XG�:�s(�G�2�!� t�:�'��(�?���1�R.���Ň�R�q(�Z��z���c+9�eZI&˒d�xKX{�n�yW��5�z�>q5�V�?+D��m_׻g���4);Ζ�a9��n��m&d�Sr�?AXf�H�?�Ɔ��U�U�SL�k��T��FK!V�ߣ+�����-6YV� �b�E�&��Cg*�Yx��)S p�J�9O��Ӓ�>���N �8���=�B�D�}z�5s��# XQ]�Y~���~�Xk$�_tH�ճ�������?�cK���l��}��f0NֹW��8���O�)���*	��m�������X�kA����h�X�W��QQ�m�~�~���ۗ�^���w�CƂ0�.�[��s'���0���ā��2�~�c�� �ҤʍK,�G<G&#�4G�y�X�{P3չ�BCkB1��A�o.��r�zn���bԅ��O�l^���p�Ś,]$����w�&="Q��0ԛuJ(���f������C��x-������yA���cǴH����x�ό�M�v�e���"toe�L���ؚ�"�T�*��; Υ�&U|Lhu_Ⱥ�D9��#��}cX{=W����<w`	��'Y�J��o�����*�,����@�&\-'E�[[m�}Cg@~��;M�L�`�N�K:��ʥ��lK�F=#���]�,��͈ `�=�^�yޠ��A�9˽ם3b��-mcޑ8��q𩑀^,�p�7�'�n,j���c"_f��eu�yJu�Leԥ��	����VC^��a#�W�BÃ�
�X�nZ+����_b�-^����4�2�;��ݓƾ���3ee�j%e�%�Q�YĻ�sr��{��p� 1QÕ���2DE]�[+�S�'[�XD9w
l/���'���m���}ԈKB�%�H��tt}|��Sv��I"�=����������;���t��y�)���57.�$�W��?G�S�����zKܮ���/L��l�����w�t�����-���$�3G�Yp�>��w�	�-6�����M׫��x��+!!c��9a7�ݐ��W;v;�T:jR��d����Bn�|nDL�q�m7}�����K��2)��x��?����U� ד4��낯oyp���'KZ�s�W���D�R{A[坝3�� j1��\� ��N�������ym.���⌋fH�q] A�b(�&pl�8�41�"�D
�s?���ǆ�N�h=`��LpnZ��M&:>՝lQAF`��[;�^5��VrftJ��`w%�.����g��7X��I��0�e��g�d�{`���2���^��?�������_]����h���g�:��m�E�QK�`�6�4.�́��z��@#���@_G HL(Td���<�8���ezH%��Q�=�(���8�P�I�<���d�jQ�N��nW��d����V~�9u��è��" #Ƈ�0g~l A�4����s:;��Qù���n����p4#�B}�͂(p��c�S0������ol� 飭d9m�T�*������`QZ�1�8�Y���E��F}��f����&�	�}p�U��o�x�G��YE�s��6�h��o����y���Ha����A�Ŀɩ�WM����1%�T�{�lp�pA~OM���=ѣ��қݵ�J^�^,�`��w� auS�lH���#�h���N��8wI��jn��dIԔ\!�=(�Xi����I���(a��>�J���G�}�;���k{XC}l;�����b����Į]�0��|b����G�tO߻�ؿW�!���$˔`Q���l�jF�f=��x�U ��r9�4���<ԩp������5g�!�uQv��ڶ�jL�ė�id]�=�"�{I,@^w� �š�:����1�G �l¿�ֻ�9�V|q���� I�98���0�Y#x��U��nxwOMx��8Q*�A�aڥ��*�xE��a�deqڏ�>����T{��ũ���לy�R�N�Z���_�����qFK�ۡ�a}��PJ�N���,��+Q["���[Ide>�l�n��>�q��f�F�ۖr���}1��q~�7:�/# A��
�bE��ܡ�)ŵtU�^y�P��ت��2܇�C4����Ԩ2��݋�j
�� O1��R�~F�!7�
�A,�!�vշգ*4iJ?��i+/��¶��~~�=�P�j�8��MN�ӊu�á��ŭ:*�5"PIZ�zpa�W|%GVDU���l�V��^RX ]�%.�VB���2��0��^�>�IE!?=m@��?�;�95B�䂚�ω�������6ҍC��o��	��U'L� cC@�����
fR�No�O0�߰;���MN�vDvE�ezZ��{P��q�l�-�1�ZK�� ��*�|�v�|oQ��-��!���^����ݚ�p�";�������g�(�C���F�5�������>+��}d�	��к�?��kb�w&�Ey���]w���zH_�|��E���z���:�l�˭j�ܓ����|e�$KYQ#�Ęa�\a��y`3ҩ����G5N�V��q�����#������Pq�,ڟn6i����� ��߈�Ra�.�̭�[u��n�'� B���E��v�Az�O���.���|Zc \�^M�__�9�/��#��q��Ru��i#�4]�Ơ���i�E=/o�����D�D�n�l+\����d��I��x*Ŏ�B�{�i�E�\"�ڿ;ҥBÈz9�<s(�C�����	/��~gZ_�cI4�~��S⑖KeB0&~�^�qw����ۆ��4ŜAdO���S�bp'�4����ΰ�o�Mr�v��t��ݸV��d�d�����vjYݰ��&�ț��3��{�w�|v���W�h9�@�(����SZW�	v�E �^��ār�}EG|�>ɜ쒰Z33Q��6��'��6�v"qU�K9��=����wL�q��P��e?;G�*W�`"�P�
�QuN���O&�%�z�h�x4�S!�B�[���m�x�E1�����ߏ�k��)~��J�{�^þ"�[���?�bR{��˟���!�a�7����*&��ԏ��+s�&���Nkb�Q����ż8aX�d"L�7j�0h�o�F��V��MI��LC���fk�䜈�o�ky~�+i�W܍�/��W����4�<�V�W4Q�g������3���h�2��d)P�X�u�S3�E��F,'�#�T�gJ�؂,��b|i���A�����