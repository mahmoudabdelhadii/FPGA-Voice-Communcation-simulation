��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��,�y�}�ǰ�=4d�H���`I"��W�`r���T:tB�T4D�m�)�	1��I�t��
��8(�8t>s)ו�."[�漆���]�~�]��;�O(1#5�-� 偙O��QZ��~rL'�x[�i,mׇp���O�I43��4d�,�H�����SN��d���3���r��m���̨T�I;uj2Y� Er�*p�Q$Gm���p�V�`�2^���,hz�<p��l�Bxt�5��s��\yq���#�@W���f:m��T�	,*�񞭋����_��㧋l�	�\�:��uGd��PǷ��N�I��_����Tuv� ���us�(H�~�{2H�:Zor�Q	#%�3ˠ!��iS��95�,?�.���/�F�i{#���Tp5����Ҥ0{%���2vpn���X�����@l����3dc�ק�3	�Ed&3�ZN O���z��s�yxӡt��v*}ԫy nj#��lc��m戭k[��5)�A#�����8�!�]�Z�s�M���t��w�!��'ÒE�rv��Ϝ�c@<U��\tq+��&|�&X1)C�����r�A~��B�&�����s�:n{p��͠R�X⺂L^��R����c���f��J^?��ܣR�O 1�rV���:��T�4���AD����˩�F�w��)Dm�O�b,�a���1$��c��7t[i2>�ޔ0,S���󧇳Ϟ�ᒨ�-��}�!6��Jyv�醊�^_�(�H�(y^����o#����X��3-�k\8�M�T�"`R�DF6ȕ� �,5�;Ҭ C�k���1\������k�t־9�}���� ���QHF��"��t�9 ?��{E_�7��!����](�S��0�q��w�9��=�i]�1�GʦȪc�W�XC�|�$��}q�6����zf(����լml�dz������*�eLD�*�,�m�]ہ6����D�Gw� �g��' A��)�m���b��ӎ���o�6ūvO��=�W�������}��	����z
��z�&�P�K#�^Qץ�_������&�)�ٺ�u#uD�	' �/|�qf�M&P)�tL�x�?�u�����ҽ�����*c"q/�\��YDl2n֢�vtX��Q������ǰ�6K�gVL��ο��Q�������-�˚e��"gb�_� L01�D��ثU�8-��Nw�@�$[�>V,���6�����=����{>G6��v�����φ+Y��	�d�A��b<�)��Gp���k�(�vWu����!5Y�N�z<V���_�T}?M�����3���[������"q�ӛ�L�&#�.~2��l�g�
*�R�Zˮ�����h1��V��Ŀ�k�}a���î�deI:VH��;r�-QeJ����f�p��߈� �׈/��	� /�eL�qq��}9�����k�#�3ęh�ڨ���-��7�m�Ǐ1�$(4�v��ˍ�HKP�K�F��8�#@W�%r1��fs
���pd߭3S�6(�L� �)��d%��'7�E��M�4cu�4����,�����N�ga��C����I����:Tڳ��pd>�s�J2���9Q��c3FP��*d����I��Cb~�I����s��D�s{�0���kH�a��j�h��5�9��&�}��Wd�_k�, Hs���V@b�q��������m���^�,G����X����똖�a�E~"g�Zل��r@�����k�sд��@�e�e��f����V��p�[���ub[��j���*iC r����ę�5����+�ea�׌�AL��?;5G��^�!l��!@�����B�佪�wb4���J�K����t8�W�ݯɶ������@�(r�.��0�@����ݷ�D�����mIXk�����q<̴d���VʒG)F��ά������8�.C�>�>v\<�<�����10����n>{�I«2�w��i�S�Z | 3�p���HY�?d:D�M��)�'�����z�L^6o
�����f�����K8�P		L�ZѤ�� 5�/�M�H�{��M�BG$��'M̔U�k�XZ���ƙ0��0���'�2��a֧6`qؐƔu�iM���f\�E��2�Ƃ��r)�L�2�:ɤ�3F}��ֈV���N��F����y���2�l�u�p#B��d�|5e��Hg���	�_�Q�YLɆ��Yi4˕bR,�p�[1��*2a%��vE݂�d�V&�
��%f��Oz�R3Gh+�@��:����Ֆ|�ױ~ ���TlGjK��q<fh��c)fg/v"��JB��X�/P;9G�Y)�+�9*���&��@ѭ�+����C?S����ќ�Ž'����!��Dκ��=�=��5<��cG��lU������lꈯ��[k���d����Zn�f}c:B>eK��T$�q�5��#-�O��vtYE���Ǥ
y V��L��j<"l�˷G��(��(6$<ܬ�����&�:�u�z�ܓ,1��X�G�^iG�y̑/�9�{��w��2՞���C���v&����L�����H5�
m��tg _-���əc���;��i~9�q��꧑�}�V�aqWKmh����V���a��D�'`��m���/1O�ٳM�r��9���	_di6p�VU$ي��j�F/���s\]��Zw��oE��GH���|�T�'n��
�\�_�n�y�����rO����7���A^�,5�TvDM��l-3�����K��Ӗ������#߼�<��$���5_�{)��n��J��x���k��X��v�z� ?�~V����A�ή5,H�颽j3Z|𻎴D�]��"H�ga��E�g�KLۋmu�B�	���*1B�v�c2���t���Y ��%��6���W��g6�A��`%��:ř�lb���waq�'�\,HT�p 0cQ�P�		s�����ƌ������&K7��6j���`z岼�^#�8f���E����zU��+���
Af#1�Y$5!=�#N	l���|��^������Q�w�_Y�D}!��:���%J�ix���o$Q� ������%4M��6�e���?jV������]�b&8����(�;�kخ���;p�)�����zl�FSCU��*��"<�~7D�O}ͪ`G����25o6�w���~�n��ֳ�F%�]�����Go��M�_HKI���@T4�#���@PV*�A��}��kX JF/w�`�Cf==Sm���*���F�膧\N�x���J_�)��� ��i�4+m����;f,�R��BI#y�:4���0.}y�
��2�2	�����j�s�l�,��U����+wg�U-�k�5CZ��}Z�R��J�T�!�@�谓�n��6�����\����?<�pJ��;�@Y���@�0xS���*0����wMNn��'��%�Ӡ�W��#��#�<i�r�;�M�E��MD�X���1%��;��l���h������������睘ӭR�-;T\�]B������t�=]�)� ��d5����}r���Mh���U.0�/a�2�մ&�f� ����%& �U��V����R��1O���ɝ<�H<�d�����<�
�����n�xſ�6y��O�`�G��t	KA����b�Q��?�و��eߝ������¢e��%�VwY+�H9���*�T���f-����4��鯘!��O~���rle�3S��y�K��܃j����K��nXJx�,��!س��r��K����f����'Ƃ���.`��]WmM�1C7_~
j1T?oy��h��Dka0 �] ����gj�t�sX)i�¯ޑVj��m0�,:f�u-�Uj�@XI�p��jt�R��e�[KS���8�=��� �x���6�f���fJX�����������@�wW�tT=e�1e� B'���=���7m���Q���gtѡH,	v��g�Z�MG|.���$�g7ک
���\�D��'�쩦�m}р`�dܕ����A�ܼ�,�?��ꥤc���#ΩUI��.)	4�u~E{���m��။
��K*Z��w��K���m��?.*K ;���ֽ���C�?���8�@��ݑ8<�dN��2�x��%��1�mD��i�R��z;̵�т�|�9z��'�Ao��KW�]	v��&P�u4�_��ɳ����	�NS�d��X�(P֞-EL	�`������և+}�a|�"q�*�	ԇ�������o⥶&�`�D@��8�эhZ6�d��<�����%��Ly�J��j����,�7�M]�=��9���Sn�%�<�f�h����݋T�q���K;5:'TDa�W$Ȳ�1x�r�.}{�Ϯ�_Aن�g��D��?W����n"�O�������$�%ɾ�KbB>���Q��E\�ww��Ȫ���s�$�E��ĵ�����-��O��;b\��	F#>����_�"�bB��m[��/�+SL�3��\q{���=C[$e�<����q�� ���?�}^r�X0����ct^H���D� ����	�� %��3�b �1�Q]����=jLNo鑂�"���2��p�~~��G��_u�μF��FKS_��+�1�{6�0��ڧ�����w$��8ۛC������m�xj"��"��)��ͥf�i��x����= =~�E67TLL�8g�k�0�jW�M)���B��s�qd�+�,R�y��4�Nu�s%e�Q�4&�GvJw�sim��l�M����q��Y���B�բ�q�R��+�פ0ƕ�j���z�� "8lf����C�춶[��Ua\J�k�Wf��H������׌� �')�7Q~z$��������e��|Kz��k\7}�v�څ}�����Y�;^$�j��C6�X��g6�!Mq�U)w5cl�V�?�Z��T'��*W�k"x�7��h���
]�d�_V�C3�G��P���NQ�t��}=:�p�4Y��C�a��_8���{f��p��՗��5T���\ij_Q$ ��7Hz&��Q#�&0�U�2�U#� ��<4:�
��1�;w�"�\�L��hf*Ȣ�*��;�j�wU�fإXfx���S*�}s�5�/�h�J6 w)c~��9������ -�k,�_�X�z�"��7����9,H�p
O-���RF��	2�|��?���*&�m�7
B�Y��bR�c�zf�J3�������
Y��r�e��a!�)YM����S�<�a>�~�ַ"�\��de:��ßU v����Kڎ���(�t�.�V�=������yS��sF����˶'�0{NYv�cp�0ꓘ7;g�d�\˫}�&�	���
���Y{ۑ�?�[� �A�k\7r4ʆq�����ǿwV◂]O��d�W����C��	"3�	s5=z�R�<����Z�ZJ��	F�e����N��|Yf�V`E�<�t�W`���Hw����F�_�7�R�C0� ����Tx���͸�v�$�_!��Ӱ�\k��BN=���q��^�\��ʯ��z)�5$3�TI�'E 2�M`'R���V���S'��(B��7��{����7O���O����(q^�w���tR�U��-�g~�p�Er�XaK���UOH_�8aճ:��Hgo�W�k�AB$t9���UC�<�} ���ʺe텄���-�7f�w�ꓡ��0H�I�3~N��<{��Fw3�_����X���%
6<� ��?�%Upĝ��
=Q	��:Nt%���,�9[���ծ8ңΌrBlW�G�&��������#��Ў�������y?���_)��1%��J�Cg�<���t\#�2+�s}��ԭL�|��U���W�F��v���������m6�0������wY1� ��{�׊0l��j������d_�d�6��@�Y��}&���h����S������69��:����%`�W*xB�Xh߅y9�r�b磰�� 0P��	��ˑ:�.q���.`q��v��J;��6����X^x���מ��·��{g����c��C�}���/Quw?�V�+�j���W��d	Ѹ�%��:�ָy�b@��,������YECς¢�:�MШ�@�jLa$1I84�|��}s�moB4�v'{k�y��m,�x}�����p�i�hC�4pݝ�y?u]����y�--�ş�,,�x`(��?>���I�`hŊ%i��O�!D�$O��z��m��?��"kL�#��\�U�vJ�����8�fƏ�#��<I�8LVѣFߒ������<)\� �ѯ��*���$�ҎA���UdP�+������LI%��ճӘ�HE0͇=�9+wo��w���"�M�:�8s6�R��T�p�HVF���Ä�r�u��9��X|�+.�ђ8O�:�m�����ڬ��D���ڶ%jIu|$'����Z���
k8��#�����-F����m9!�K�q����uku�.��T�gĖ��?FY�(�(|vֺ/���|�K܆)_&*,��\K� ��cˡy���$�r�liQ oc�t�r����r�rGʞ7
�(��+_�:%�.YE���TW=��T�$��+��Jg~���A������t�*���-��lЂ8 �{���g%�f����cY[g̪&�H���f_����p!�k-�ϟ�	��K�����Ϻ�`<(A�B���V=Dw6���38��f��f���:)_ھ�,��A�J���@7�/���i�w�����l�+#����R֩��Gdg�X�c+��	G�V0U���#�NwtyOHb����%+�s�4=.�/XN%�K ���j|Yo9��B\#�֨7��uIS@T9��K�溇�`��;�r��֝�4�s[�	D%�E��Ŗ�8LO3ψ^Vf�1�i�Șk
 jO�zS	}N=���~���KH��Y`��u҂V:�_�]�s%��n��z?8]��Ƭ��m%~b�MΊM�Pi�k�OF�5�꠼7�J�����˪�3�4.��m�y��g��7�ab�O �p�����������]���2?�=.��I5�5/-c�'��G��c�/ �&�Jy� v�e����䋯�i�>RV�j����S�W������iD�o�&=��}M����9�T���>Q����J��i�=�"�^��4P��9Z�r�p�332(QAKbcaі�r����JA�$M�9��9�?��7�|3�fpfWg��;���z����rBt62G��,��7��8���p�� @n�>�s��
x���od�"� <J�od�e�O�o�<�Z:B��<�pkw��awok��}}�eq]�<g�{��'�fݟ�p��O��ö���|����N�/^V�͇��ld��w�gDl����5��8�x��Z?cy�㺲�eU��[�K���x`��Lvb4t��/�>��lcA�m��V�9I���e��5�S�K:�ō�$���c�Ut}�w���; �e�.�z�fT���M&h;��E{�v�z�b�[sL0u�hĤ���-3AV|��8����ۻx�Ǵ����#~�N .�Kƀ\��L��u��q)���x �l�)B�1ޅ�>�H	{7:o��_���N�'�-��Y:Q�+�X^�h�|���wDY=p���OAd�����j�.�?��	���Z�3�L?0V*?)�'?J�����61�bK��+�s�Z>�ZL^��]k��rL��4���f�[v� E/Ox�OS|� ]��lGX���������E<���/�޳��S0a��3#3;O�`O/�O�̯_�hr�-�U�eW��"h�JtK5�������v�@K�><�fZ� ȝ�T���}�2]�<ֲך(�|A�=�S~�12��7z��R�~�t����g��	��B*n�J�'U=D���II:�uQ�s�Q�������!)Z)D���?rB��'�n��'����v�@���t�O���;��C[I���Q+r��5,��HĬ+j���	�����)~�S��4H���8�Ƃ'Pj�2R:v`Uee�E� �#�I"��1�UBkwOӓk��C"����ef*�@N$��Rm�b��,��x���w���ɷ��n\R���J27~3�?
7�Q9��A���Y����iY$5M/�Y�M���-o������5u&r:+����x��W_����܁rL�l�M4��&��[�h4���M�YYM(-}�������]}�L��)z2,T�[�O^��5`T����`�㳵)1YA��d���˞qd�^�3�1�t�����=9�UJq]��
��l���=Z\��si��kg�-��DrS�4hp���|��V�X,B����M}�G��d`�
��Q��X�>���}���n[�#�V�}Սr� ]�z��[�������X��IЄ��C��P�7H.���P/������o���l�9k��qL#��B?
`f\XtC�sԓ*�)�O.h+	�Y�����X5�x�y��#epi �;$f�#3�+�d��<�"�����)��"t�O�/��k��r�murnBrM8�!��*Ys���C��P���*F�{f �Ĕ�1�b(��[>�fg#{��Y/<�
X�ˮ�nq�$�[�/G��F!��h};1�׼)h	�9��i~!T�"�>"9g��'�$S��k2KK���?*�w�C��v���-�cҞ�w��%=�����|(e ����z*����$~�"b��ۯ�G����C���M�,50�t��
�t�r|(��~=M8�S�i:x�^�0]���9��/�2�7G"��8�O�L��A@V�Z��,���p�ėj�Kȵ��5����R'���~C@���E��5�p_�Nم�D��H��ս�C�{v�p4V+�G<�,����!�4P\qyj�-7�����$�Z�����[�7S�|I�.q��t�+���TT��}Y��|��8~��Ʌ�a��I��J�7��s��)��~\N��"d쯐�͸�~�E*�3�c}f٢Ή1�o��N��cC�j�0I�g��ʛ������ܼt�pᵀQؚ2eH�!n�w��Y�����F��1�[⭾t'��Z��.(w��@n�����^|���z������m̃���!��𦇦��Ao��
�y%���l%||��;�<[�\���I����Q���w0�w�!p�=b*%�O�lO(�MK� ���%B{-޹���k��^5DN~``�m(N�-��A�9�%�K��5���]X&�ۊ���+Єs+�=ͦ� ���ᮜ04�Y�F6�g^�v�,�v��^q��s
�,� /��A~p��uz�?�NQv��T���{lp*�Җ������%��G�B&\�AF����`����I���~>eȍ���r~�{�/3S䥿�aq���'W�s�c�E�l�*��gU}!���^�k��� z��1�;+�"�4ȷ��<��:m`�l��O�^^r�L+w�k2Dw���&�!=�S�1Z���8JפF1'�H��i�M��( }|!X��}��\�)ׇu_�/��壡�Jj�/*�vu3���J�mY�4�a�{ �f���'Ã�ߝ��8�	#�
>9j0�$�轣b%�C)��j(�y:��e��eH]��Fo�Ҏ	��?LG�@IlZ��b��\�����ݪ�C�������M���+����k������g�˃�Z�
�b�=(�kX�k�\��܋'��P�KrU�5������&"˒6c�S&�P�$�R�0�c;[��&�H���(�f���a�/�c�Aki�X݌Dc���u�lT��"Q=Wf��O�Ty���V�hY��0q6ʡ�8��*�Evg��U9$�Z�/K��{�#���;���un��������՞�w�,Ʈ�w�,�N�:���g��P�D��}j�#���0뤣����6��KB>>��sz8�Z�n$B�9��������:�ŵ�ܖ�_
s:ʅ��DjT-�c����#3�@�E0�T�6��~�@����'|/ 3�X<?��[R*�����*��:�\�Ȑx�`�����}4|圱�F��O�
�ʦ�?��8C���U������ޅjv��d� dy{{���k��\	>�f�XcǗ���F�3�
���mP��$�}��vy.E��=�{�:��{-�/� ��`�}��0�Z��g�Db%�r�U z���n޵!m�.,-�P����$���Hjq�V�2�"eb+��Pj��t+��C^��p3l!V��$R������c��,!�{=zy����za"]��u� ��g4_u��^���I�Zń�i|O�Ҟ��C�+�O[�gJ���uk�P�7�إ�� 0��ײ{� &���I�A�"�?Wf��Y������9��yg�'5�i��h�B�����P:v���:���X�Ȟc��gXX({�c$�"������i'0�mZ�(k8z���$�<ʈs��ST����1u��X`�]�B����4n3e4<�e�:�~Zuha��o>?��~��%��~�h��;	���j�c�d�4��͛Τ�����_�$������!~�����';�M��Y�&�P�#��_-��i������U7AG�X�G�׮/$\kCD�X��Apo.
9��9F���a�_��H���s.-.�:����
��/̈́O���9s�,�?s�r,�T_ˠ�54l�ta+7�ʢHH���8���5��>^š���MXڍ�*������o�����e�G(����g�Vn���&�i"Y۪���ʖ��<��)n!iT$�|��61<m����LـY,b������t�O_w(�S<D9��bb���>�oL%be��n1�s�ߺA��Tls½H� BIO� �����#p�f���N��?�50���-:�\�∻R��R�#Bk="�� ���F,x�Ĳx�Q4�_s4w���b$%���w�	�;C��J�Ҵ��*	�[=6"���|h�S��H-�*� �k�����E��O�,,��ˉ���n���Ɇ^DcȤ YJݤ��J��f,�/6@Zn�<�,���D%���w�<K���j��c�������[�����>N�^�`1��j���]�y����[t�v7�~�E��f\g�δ��ӥP�I���C���_ �o�M�R�B�EE�zn���ҁP�Z8���o˒�.>r ��X��XoMp� p��b �U�Q_�	��MD��m��&a�Ϗ�}���RN�p޶�m߶�_�J���3�ő�n�D�J����	&ϬH�kܾ��̴>H�A������ҡId�%o���A�c%�5I �5��aa�8!�Ȓ0`�?˞v;���~����E���YHN}�I�"}W�������E��cUU��U�h;�����8�%{��N�=���Q$�����]����� {�P՚�{�i��2�hx&�SQ��Ml)tw��V ����@B��U1;q��� 3�p(��̷�ڧ���ה��m$�h�4�QƠ�(���t�#?�o��"���)cb��/�|�S�"K�2�Է���w���c���C�P�j�ި�S�X��nf|ȃM�=�/�Y��2���:������׭������׼&�I�T�h,j�iT��*���^{�`#������F�>��
,�SLO�A^��;�ڿ�p� ��A�eWu"��2��Ks�Hk��k�И�@�UT	��a��B��&�����A��#����(�Lz�D�	�Lf
��;h!�T�%Iɍ�����E���ؖ����N@ &H�Iz"����Y�+�
�nkI�z��|��@�]��Dv���0J�f3:�A�%rm,d�Pk�yy.�^�"�)�-!9G������lUh��%����Fx}eH������-��T�6]���F<�u�g���o��	���-G���s�d�bt�)ߤ�s�M�<eH@O^i�灈�dup�y���n2'页/��$cI2��V A�V_�iu#Xt��H���/m�),8ײ���hp�8��yg��&�
m��OZ��wrFm��;��z�}�N�{�E3X5oW��B�X�=;K�٪ߧXyo�!A�F�ԄF�g�����-�x&�L�Y!CNz��D����ϱ o@<k��6�ʢV�Ӎ�L�_����@%�a�LۮrJskk�@e�4IJ���{
xx������{�(r7|W>��l(s-�m��n-ğ�6�k��~�V_G_.V\B���$�.�;w���#4��<H���g?�$��
j�,��9�'��Rlrm�l�$J�/)����'H+o�8�E3�
6lN�ӃOϿJ��k����]�̠�ψ-����wZSM�)�(X��F��"CǍ����`�rh���%xK��g@!^p�11Q�6�J�h��U ���h6[qڼF ��=�-���%?�0ϗ=tk��_t�t/��:6�n���󒎪��KE�M�9H��?`iu�jA��qk��SZ���=����`����Px!�O�d|�*_�gh{�əx��V�-&\@}L��x��+�e����t
i=�G:^�*�����sJ�0ʿ��s0ҝ�O�E4o�`ȃ,^�ˤ�N�P����V��9���؈x�E��dP>AsOe���t%��2[��3{#�	����N��� R����Fq�k��V�E�x��@�V�2�z���z�aO�YĄ
��'+w���?U�b�7����i�Gͳa��|�҆��%�O��_� ls�d�+��TR<ʆ�SVI��+��;Y2(-xf�!\Q��N�V3���5�5!˶���i��5� �P_��@@�P�E���Ԗ8x$�M��0�:�3S>����m�b^����,$$��1�W��,�E�2�x}ۗg���t�n/�~<*���g�P���
5oH
�19ʤ�������Q�Z�\�*�t�|K����r<(�D[��ZE� �)�S�������CX��p�}�$ta��$�� |��t~-WP���'q�d��'�8�Ư
�\g��Hc����|l�A&ݕ��d�G>|bơ$�R�>듿}h��BRs��?]ӂ�?[�j>�?~����S/g��(t��������*�������P��~�2��j4jݯ��Ӈl��B�ph2c�朦��`�������f5���2<J�]��nt�A�҄�M<	�Fj�mF�*��uKb) ;#Ͳ-�h<1�ly�2l����?�N�7>Q��
4Dw�33KG!2��>�':a�W��j�u��4���>��P�pf�&��t�f@f��ix$�� 3H\`�4P�@��,O5�X��@̜X���`�