��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��,�y�}�ǰ�=4d�H���`I"��W�`r���T:tB�T4D�m�)�	1��I�t��
��8(�8t>s)ו�."[�漆���]�~�]��;�O(1#5�-� 偙O��QZ��~rL'�x[�i,mׇp���O�I43��4d�,�H�����SN��d���3���r��m���̨T�I;uj2Y� Er�*p�Q$Gm���p�V�`�2^���,hz�<p��l�Bxt�5��s��\yq���#�@W���f:m��T�	,*�񞭋����_��㧋l�	�\�:��uGd��PǷ��N�I��_����Tuv� ���us�(H�~�{2H�:Zor�Q	#%�3ˠ!��iS��95�,?�.���/�F�i{#���Tp5����Ҥ0{%���2vpn���X�����@l����3dc�ק�3	�Ed&3�ZN O���z��s�yxӡt��v*}ԫy nj#��lc��m戭k[��5)�A#�����8�!�]�Z�s�M���t��w�!��'ÒE�rv��Ϝ�c@<U��\tq+��&|�&X1)C�����r�A~��B�&�����s�:n{p��͠R�X⺂L^��R����c���f��J^?��ܣR�O 1�rV���:��T�4���AD����˩�F�w��)Dm�O�b,�a���1$��c��7t[i2>�ޔ0,S���󧇳Ϟ�ᒨ�-��}�!6��Jyv�醊�^_�(�H�(y^����o#����X��3-�k\8�M�T�"`R�DF6ȕ� �,5�;Ҭ C�k���1\������k�t־9�}���� ���QHF��"��t�9 ?��{E_�7��!����](�S��0�q��w�9��=�i]�1�GʦȪc�W�XC�|�$��}q�6����zf(����լml�dz������*�eLD�*�,�m�]ہ6����D�Gw� �g��' A��)�m���b��ӎ���o�6ūvO��=�W�������}��	����z
��z�&�P�K���Fn�kU,{��:Ծc��%(h�=u�ݦ%��t�|+ǆB�������0�yȒG�좩�����h�g��M�����!v�+���#,F��iS�5~i�� �ؒ`.�|NT0h>�~���M/%{�mh[����<ljd���P�Тi����F�Ϋ���g��j̆g^�k��k����A�s�ہ?�%�C��;xd�ǘ���.!A=K�,K�9�>�4�4��[I�בN�^�Ha"=	 SLA"����Γ��M._��w�5��h}���l��7:���|��	�wS���=����XZ�^߼�B[,EJ��|q¶(�"�Ui�x2a2��H�A����-�V]��4����X�3?���Ev~"k��æ�c$�L���S�ӥ-E���ݺլ�!�}��JGD�����	[��ٵ�� �2�M�"A�6�����/Rh��bg����
������DQT&U��u����1�
�:�;m�b�V��bk�^Mmң��+�X�*�[:�`�\��x#��S�+M.6�㿳$z},�
��So�}X"�a�S�Vy;,t:�����# W\&6�TIy�~�{�9�
Ϻu96�)�t��^�孼E��X����l�_J��<��#�G��t;��>6�T�S4�P�{���X$���MN\���,Re���D!z�gx�@�}:��4/Üp��vأɯF�����h�3J`K�Ft�j�Q)��{��ޠ��)z���oe�u�P���.���XXÊ�T.��4<�*X �=�]�?@��(Ӌ9�Z�~����g���~������7Ap[hD�N�+z-0QlC"\s�5&H��Y!�`Fb;���DmUө�h�:�(�~��?	���bEЄ��_�P:^�ܳ�βn蜫$�����n���H� H\��cڀ(�߁���c�'Ht�1-!9�L�D�|��~�E��ń
(z��������~��z|Rs-��qs3��)`Y;ȝ�������?���@���v�q����,_d�ڳ�8/�&*���ӱq�Gӷ"��[��He�U��w��(x��B�C�íkg�~>�N�WwإX�1(M�-��C"<vTO�b��RF�FJDw+�FV�[B�Lӛ��e7t�P҈*/2ט��o�9P��[lg�,L��a#�P2��|�יT���C�Y�c��y��Z�P`����+	4�IAv�*_�����<̽]�U�(���OZa~ilEH<���W��\�9`9��s�䣇ـA:e�3�'exh�q������mEG�D"�!Gv���-c�x�f���z�&��l-r�m#�����Y�C���@Ch`�V�� ������t"gF����X#�-�	�&y�b)�'�4n���s�'f�F�:���?3D�i�Æ�j�O����?��$�����u����,��t���(B3�6R������Z6pd��EBZșc��i����5:�9*��t���|/pW�T�%�4�AM����ɜ��)D���>QA���!�*�Mx-&U�	k�[d�
4����g�wk�`ߚB@�K>'����4��A��V`r�J��E��y�B�Q3��t�
�Q���t]��y������Ӎ�u��}�}j�(�b�z0Z���M��^3�k�:�3�}0��<z����N��n@�ʆ���A�
��NsV�{_��zFy皁Vfځ�D��H0��`B�p�d��ֆ�B/�q�nWM'մ�����҂��D��!΁��J���d^~TEI��I*y;�ݻ�(8e�ݻ��t�/� ' |p~��22K^�hc��X�*W�O�v�s��c�|k>�)�������pJ\A�S��?����?��v�����w�@�R
{˓����2�E����Zɍ=��m��XTz�gw
E�t&���* �o��+�b��f�˵���lۤvR�ck%P
\'�@W׶�k�ٷuor��� ��7^��GG� J���SH�ᛇ'a��r���4Rq��MΉ�#d*)��5������~�L��
fKo�n6��f������ �
�>�K�,jw1x)�E*t�&2�,�O�w9z�s0d7���႘.�1~z��Rte[ʄ~M��Hد�}��Ho�j���Y��a�X��	�H&3�w�֑�C�7NȞ�@��	jn <VW�[�K�-�[pμxd����#��,	��.�я�iii]����*�R/x�ũ�����P8���O�j
U*���j@a�Bq��G�pb;��z1�Q��s�^/O)��]q����:�� �trj�|�j4{���7n|;�Zhmn�Q��������*&⁨��&��Ycu��RV���9,dD�S�V�5������ذ50�F���k]f��u�G 傤)�wf5�gݷ!���L�$bD&%}=�ξ�&�t�?��Y�u3��T:s�t�� Lk�뵷F6��h����-�CG2��g��@gn��;Ȩt-������ ���c�v��}*��br���,F����ք!눇�7v��F��E͝�����M�Tˤ��H���@4�K�x��]����p�y~$�yDF�NAe}�0:�9
��*k�Sd���s�#�D�K��?��kR�rCaWm.�=�^���m���{$�iS�?���+���!� �v�~ǫGݻ6?t*Ik7T�_�i�������"<��WwA��ܶs��e�P;ʜb��X&��?�#Mb��ӍM��"�Ou��%���c=�=忶���a����*#\Z|T�=�O���A���H��Y6Qp 0���c� 8��@f�ң
pnO�+��{��	��`L��ᇵ���(/�J�c�$yĠ_���.���d����(o�2�6�3>��~���JGG3#0�VF�,�I���@vaQ���L7s�x8�*�QK8���������z�57��6��K����D��=�0HG�>4�q����1��H
w��m�9�� �w��0u�$�п����g����!�^���՛�+qx(o��!�<��c�D��D�^3*٧f���q��`�/���]��}*���E���ѷ۱c)U	.��+>��LTB`��B*va�b�Ŭ��C��Ŵ�'��G���
n@O�$P��m�Z���9G}��@O�|������j�?��?�y#��4/Ǚ����	ybA
Z;c�;��^���LVἰ�Ej�awwǕ`�S��-��8�5~M4��f	j&�̔?�zA�zj�n�b�<nN�BXu1�=�C?T��³�ҡI.�|P�MVb1٠۲�������Z�~��gػ"ņT�%��,��P��qRo���{d�Ot}��������!S�Q��ֽchٸuO"�8=����k� ` tj%� �4���e_��0�_h,�`������L2�4���ٙ��X�a��&��)\��t����y(B���q�P�hk�R��.Ɇ$��Ά��H"���������oƢ@�����J-���mM�c�	x�A����<�MGr�TS���H���+f�V�
_9�
�˜ۣ/���Rh�k)	�xM�N�:sˈ���jQ��/��im�P�D���Í�N�4>�����1@��D9�K���pDq���[3�",����p��?\^}��%T��,�]D,�����
{�� x�=P;�k�"�fI��%���B��g�QJ4Axh6􇻰�afO-�7 �4��Ч���u}�h���h�P�K�$�p`����UQ�/g�w{�1��b�Y�V��B�·ˋ)Ē�#�YD�/�[1*]ʂ0�0���:ޗ3q��81�o�U+w*�E�0	u�d�1J�.�c�jX}#�ٌg#e�m��~N�xV�2�#o�?�	2)s������҆y&�HG�[
F���C�2_v�j�l
��#N�TXJxNs��8T�x���r�0؈�N���XY�@@W~��	_�m �#���䱜zo*�A�8bDy�`�ug@�n�Ǒ���Z F�%�]wS�1e������E���X`{�x �p�u/������]C7)�]�m��2[1�A���45ﱌ�p�K�$^�2q'i��l%~�%}?�Kt�|���_p],�����Ѧ�	S��>�|vM`JG��P�Lv�&ը)F\c��s3�$mcά���qe>lF��}jK1JMH"��-��==�z"�*��NQzf����C�N���b� ו >�b)S�g�WyQ�K���x`[ޕ}v���dSI���g)���"ځ�'p���=�5�̼'
� ��pϏȇ�qɵ�2�����~rP"��.�����W���~�r1� �0��#�C5��*Of-��M6)�{l<~]�# �zw���\���N���u��JCI�P���v쌜����Dm�y�\۷"�O�:�R���*��Le(A��x�h��ଝ*��rǮ.X!i�r���G�����q�3P���@3s�	�,�w��i����?�O�W$�"���ޕ1�0X���?���򄊖���J�CWU!��n��d�j˒~��R�K{@4��MMy�0�!�J��r|74Π ���Q�cV��#^K�IC|`#�U����rL*ȝ��ۼ�A��M�Ll�_"l(���ӭ��B��T���͊ %�>��n�=��Xb�a�lN��2���G��^��L�Кn�j�c�G�%cj�"#GYU-a�4�