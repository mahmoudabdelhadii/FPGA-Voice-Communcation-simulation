��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��,�y�}�ǰ�=4d�H���`I"��W�`r���T:tB�T4D�m�)�	1��I�t��
��8(�8t>s)ו�."[�漆���]�~�]��;�O(1#5�-� 偙O��QZ��~rL'�x[�i,mׇp���O�I43��4d�,�H�����SN��d���3���r��m���̨T�I;uj2Y� Er�*p�Q$Gm���p�V�`�2^���,hz�<p��l�Bxt�5��s��\yq���#�@W���f:m��T�	,*�񞭋����_��㧋l�	�\�:��uGd��PǷ��N�I��_����Tuv� ���us�(H�~�{2H�:Zor�Q	#%�3ˠ!��iS��95�,?�.���/�F�i{#���Tp5����Ҥ0{%���2vpn���X�����@l����3dc�ק�3	�Ed&3�ZN O���z��s�yxӡt��v*}ԫy nj#��lc��m戭k[��5)�A#�����8�!�]�Z�s�M���t��w�!��'ÒE�rv��Ϝ�c@<U��\tq+��&|�&X1)C�����r�A~��B�&�����s�:n{p��͠R�X⺂L^��R����c���f��J^?��ܣR�O 1�rV���:��T�4���AD����˩�F�w��)Dm�O�b,�a���1$��c��7t[i2>�ޔ0,S���󧇳Ϟ�ᒨ�-��}�!6��Jyv�醊�^_�(�H�(y^����o#����X��3-�k\8�M�T�"`R�DF6ȕ� �,5�;Ҭ C�k���1\������k�t־9�}���� ���QHF��"��t�9 ?��{E_�7��!����](�S��0�q��w�9��=�i]�1�GʦȪc�W�XC�|�$��}q�6����zf(����լml�dz������*�eLD�*�,�m�]ہ6����D�Gw� �g��' A���FX��\өܹ&�6�h�Ð�$�(+��埧��= Eza ��찠pr[�c&��nP��x�2�TK�M�V���3Y4vIR\������ɭ�1՟?4�_y�y+����ƄJMm����@����m�����c�t�����:ud�Q�����T4���QxBŎ��\o���t�*Z�$�*7<�t~eP/`lfhg��6��[nn��#<����n�D:� ����4��1��B�ҀΫ{��5��.�%�~���R6�_���Kؑ�<2��{,���!���O�Ǩ���� �U�n�`�1�C_�I���!s4��~X ���+��C+���XǄ���E}\g��٤b^>8�ݭ{�]�*{�N������~I����11�|hCk���K��~�x!��� EV�R�p���q�/����# YԢP�JAnS�aA��_���R.r�ʗ�)���
ʥ�8�[�w���'�t���u���z���7�T/���^-!bO��XDQ�(]�ax] �5�HTh���h���}:Oބ2���َ���IC�g5���Jg`�{׳�ʇ͆/��S�̇�chg]�quM;��ڑ�y@�94��CCL��弢yP��^? �3/\�~�`}�b#�yۺ5�r�4!~��:�t>�`H����J�[N�-�"�������]N������H~�"���w�cP	&�}8�1E>��FQ�@+���� �Qϱ��Tg�ϸ���)I$�	4���ʓ!aj�A#&�\���HT������W��ͅ�k�ˆ��p7˒t�TG��[n~D�s�Li�ƕث�o
p*�������@��}�-U
�ьr����zq����:[+��vF�ܔ�@���4�)79UP-XΕ��5��??��J�ޝ1����<V"��,�u\��93d���EO���7`���xm����*��cda��-/�ο�tw��M����l�>'��o�ո���<&�x���I��~��x$H���((a�\ٙ&�X�1�H���U����,.���<"�ڵz�R}���,|@%}Y�ä��Nɡ�l�'0���Ҷ?�;H6����D�Q���d��E��F�w�Pw�8f2gP¾�������
>M&� �Ȟ�i�S����)%%-�j�"�Ҵ��:?����_w���:�������ɝ��+�*ZeSȔ�ǟ�6�ÇyC=O-��nh2}D�*s�gc��C/\�HQ��6�/�"#Ɩ�Z4��x����zC�ȳR�R��h�w��&Z�GRz�Y[�d�V@����h�w�.��l�֞9�^�K�`<����' �ҫ�s$;�
���������{�}�8b#R���3xW�)��!�����!�E��3�h)�r�� �e��Y�7�����}��R}��cSV$��� ��ge�I�@$�Q��&Zc)���1�a*U�6�<�RR}8�{���&8��[�������QgP��y�<<�b��%�rP�{~Q��GV�5��1gLx�i���q������h (:��(-�,�G�2��}����[f��a���;3=��9������y'S�XPZq((FS��Ep�íCf��&iͯЀ���m�<�fu��j�\�B��*V4j�/��7)6J<ڱJ����=�EM���Pw>��Dq��tVw�u@����Jh~���C���0T�Y^�BV��pa%��褶M����b2-~�o��"��:�}�4/�i9~�}����Iq0��~�ޢ�e~��՝ຖZN&��d�֘���QiKtŷT.�
�wҍ�B�(�5C� ���<ɴ H��B��6bjH�k��`��{�	6��w�.ǻ1�i�AAU���s�}�?	��u")�v$�Xz4���b���о:WՇXu"k�E���N��r�(T�'	��sY��5��g(pI��4sJN:���d��n��䗍����?�b�;��Y��r�wk@Z��c�tD�����G���FLn����˹���=��Y��s���M�����Qs��nI����H;�I'kt+e~�g��f�62���g�/xb��ݟ2�8V�ZԀ��h�Ȃ!2�ʝ�y�pW֗1/�fz�a��͞���lU���B���;罰�%��2���V��j��,���Q<��6t�c��[t�� :����֊��#v����������V�d7�,*�����,�	���4g6kq�]
sX��F�ҿ������?��<m�SM|;����3ʦ��Ҽ	���� ^��Ax�V�Q�]O�>�9<���"MȰ��M����2���6?ߏ�6?br��{�QC9�� c�	M�T�0+ɘKkc�E�i��S�7]β�r�������Pĥ�f�Z�`�����.��[އ�]��ɉ�P��/>y؍�#�Y`�v\�rz�bdvRG��"U�X�xz�k<���J+��uZ����J+Z�d�7�|�*��Tm����ђ�ʽv{�t��q`?RI�p��S[��HjH��F�e04��
�Цf�F��e�ؑ)�h��`H�ʈ��׹����2����A������|��+�+=�^lax頄�w,݆u.k�-���f�����ӂ��E�Y�@�;���6X��n2n�'<�L�+�F6|��=��BS���n/ ����v��Z`W�3���5�/(�Nt"������tY\�a�_ik�1��