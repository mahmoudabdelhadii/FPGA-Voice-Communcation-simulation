-- (C) 2001-2016 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
ZnR1fGjTwk2vyNlWGlYwmv0UuD5MzOvYbqXLMZjzuMm6YOlmfF6OdQywmgEyGMeR2JblYiHWw4Vv
PLynxDj7MK+q70ptSLLNn4s9nGpRtaB94SKmoFHnrTY/ExJnaMbUAlgPyl8FPvCh9DcykR7zFXyA
B0gjsPSFXVQn7YUSSg9kQNRd/YaN6sIioW+x7YjrRW6s1nQvNpAWBTJfE7+Z+fOHmJ7U14ib4P1V
rXqitV4Jxz/7Oz2F7VGm+f829JqDuWVR8DD9e5XwElxlogq5q5zAdcYPWSkw+Q52Wd2w+46JQZo4
+W1jciQgjlb1cm+ZjUxgR7aU9WmUSxn60AtNFQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 9392)
`protect data_block
kG+hUuVeVZyoEpKRA8bOklRgHm59XzMl3S0DESUTPmXoBPUk2zBmnThBzeE+gcuPA/FiskKTqitO
3kFKRLSrCVW8fh4Y9UnH2z18B676Kuh/VF5sT0bFtXO0AaUR6d8i/dI5ZU2leyUq58dWFieSe7W1
K6R9cU8P2EiC3aiQLPr35rF0o4rkScscLb2CssN/bjTdRUtI2Zf2oklLSL+a1WXIzhFYChML63S0
ggtuROlT6S5TgwGVUFoPDnobok4b1PxgrYeS3Rbq0Dd+91VmXflnjDI32rgKvgxX7r+rwCq/ddPS
Ok1ZMQvHVfXsdkP0LCMQwH2SGz/tXLDMr8OK6t02v8M59gSv/W63v4nSIHOjdwC+zeDvAs783uf0
XCIpSBISZ5cLpWD3uFOR/ngD3oIQieB5ppbQaWgTNB/FPDAWbby/IRNiSbWV8nYx4Ifqdyl/D72U
ZkF6i1AeLaKTvSxJ12jOm0TufFHQbr8D0fxkMB4pOivnNY0itTJQhoqHUUHAXBJlK5+/jP7DAk/D
3wCEVA22Tfx1V4AC0cc5JMCFaNhZocSTciA5AOolhsHN3L1jyrSr60BtH4iOa6q+Rg7MLN4tbbK0
Wo8pHUKq/FyY//N1LLHZaTb6WE3tw0o7iVJbgMNi8cw4Il5LEuuwnYfb+MsIAKrX9J2QNi3DHOy3
mF2lQXZnjzGqJFn+kGfVcLa9vazDGe+8DCP8vXhvIDNq/uAc1/t1X+FLs6PGCBz4F1M0oO9+TyYb
LUYB7vl2pySf0NssieMKuR4/e0SWiDrjX5tXfv+qfbsX6+CcEeb+g/+HXVr60Krgv168cC6YYu6Q
MF/ZzG5QP38IPXfuerlUGvOycSzrBdk9KiLmDRzyrxg8OyVhyoEGvj5dsoiLirhLnVti9VF/J9UG
ljsjHQhQlEG/sxOVWXHefO4+RoMJtfhyfjzPoxcEXbRpBq01oQsNqkFvt0KQLy0S5Hgbdxhvr40p
607cYf/+nzOOtRa09lcNDLEVVWUK4Gx6KWGLK5XxkJ7eoGrpKGf9xK7LrJrK+g7E4m26xtmS8FWh
xEm/9HeYe7vbtCpcgxyADI4A6P8UK4h+rex3mVjr/pei0aMgaERYtA/PifM7f+nmHbjhmz3ReOJq
Q8xGJ69iI9etDfSGteKCXh4J7Rkbwu3HFzRLhu+u8hDO3NvREw8/ukjEI/AFUHdEU9M7B1nLV3cU
NgDoOeZ1OVwtW1Jim2EgwIiP+LuQyPvOnqXJS8IDH1Z9SZZadXMKyqZ2dvsp/q8CcFqVI66ZvWb7
6gyHHeqAEDkjhAZY4hS/q1zI6OTQdJ2+YF4bvn4ZhMKPjzgYsD8SByiv1+jw1ubBtaeZH19PzXR7
Dn8EHj3lsOW6gIjj4xDrYDdp+2/JR74pjYm0Xr5tQ2YpqLuMuI/ueIeaPXNNS+wmClFzAC+YXX8L
811JukjCiXDD1P1sDvSeXBmY7/+v+l37MauVk1o0TyoXZ3dvSwZmBKU6X86d1u074IijTb7yrJYh
vpwTFzJN1UQP4NEzHCd1ZVjM+XgQHC6+CF4GWwy2MGBZrQP+urWEk4+y7ePK1hsiR6GdM8JADkfJ
Lr7D68MnmEGnygKLfALLMGTW3WiTG0P3Rm24Osx6wgCSt/0Wo0Mdx6MUZA11zdvXk65gd8p3a+T4
u9ayGY+5n/m7TxlwJeNHKXDNPz3/ym0Y4sq1CO0qHA+Q9H932IVN9YBOov/KW04u/4A9Bl/cdSms
ET0wJkWZSawLBQawg/esJ2NbwKNBkS7ZU+Mn8D3hvIYVC2wTxWUh2WzWvHO37kW1oKYNPSCscCsM
ylvP/alPus2WOT1JmH53qGHKe+7tN/yxnaIkQ3VJXDn5kKJoZ1yN9rbbDtW5Y2F8HBZRgzYZe8FX
wVIgeeCNwBVdcGjT8t6VfLrJfeW2mAnZorYQm9JThVUdoDNh8tS1gvB7RQYHU7y+qb2ylT33LZ5N
/e70BCZIPWW2ieHFU0r+E/6j8j03IBJ2OfyRCuPpepzmSid+AD5aYFXgN0KDIuUD0sm+EtM9O9IG
ldVEx5Qu+0xRHYsdZYTINWB4Hd65oy+Hk/Hqc2uOaHhuwd8GkxpHq20EV0fE8Q9NQx8F0DpGwQqD
sFA6XyddhN3WBUlnkyb6XRIo+qbvZYFZIvi37nh4ntzvcAkrhg4U2TipwqRFsqpKO7VN4ls8zDY4
c1HOHEmhmPv/CHBiHeNezFHlXlfRR+UGzA83ncz2MkpZQE9yO5wUN/AHOOokI/aqcqnkGTxbJP/8
mjJJCeaf5e1eHUDM7ZN0tQAISqJOP5j6MLc6sitYglV2h18Tmi5EkF/mJhE/RKRmrJ20MGeqdGk7
YjGKFqbkOGy+s9vop+EnwJAAzpqjdoYypcn7F64Gv3zZ8OJEc/cQUO2lqW4Zr6Pb8U2tIgDSLgnE
2RcVZeMWQw1+5dIpsNSiQtAzV5Q5xqkFJ/pie54P/wj2AlNehsnsPGqatO7GVUVvRV1zdQIvTM/o
Ku7lVd0l0yHPIK3xWAYTvMbXffO0XOFq2IB6IRYot59GRO1nUi4pNfodlx2KjcJb23n03LYFFI9Z
ZkRgqVJ3o89iZtOrMT5BQQ9WZ8Zss55Bvkr8EF1pMAp4e2riZJw1JZjauTBWxiKGIfhYdbr3Yqp0
PoXw0HZFmFFz+Qn1WiXq9sE2hpKffOeQju+ttpDAApH4aMgO9GbOBdJ18pMGe4wgHBTksYAUgdPk
1nH7KwiD+d/wlzV3uki0bqBFxz3tR7poFRFfSdlvP8ml9Sb3jWBYrtWN/uZU0SYA+sx7w/XSbbZe
Pi9O90Z7WjlVfJt2cdNLrcFQe9Sw4qyl273rug4MPcJx3gbtgufGVDFdo6F5TVchXMgmFAJdRDnk
nxtZ8/I/M103V46/ZTkR0OUsyzKNRbBFdiHg6zjuaUbNrzUNKUFjOjdQ5FwcMsGYQH8QEdcvQ5zb
JXK8YK6FxO/6lWja4P4cEJRTtuRLWgXtwx+TTJE3nnd1neiR8+6aogNxsNKDxMgtAcxNydosGDDp
ZUDUMqHS0Rb04/JfLQW/WGxFteACUzyiP3GGpUO58LzoeI8MmKPfe52RCaOChoX8tcDZgp5Ohlf2
n7SJHvfvkTox/Uvg6Ob1nxQJRimmGv7VW7IZy8D9aDAYfv2DHkaagiqaRzJna5Lx+Xm2eB0GVdhP
OpvdOIQUlE2jAjwcSY8x1aRUvAJYjYeNhkuZ7q3N7eNG6sja+6dOcnQcMIWQrpiapLXJBM31aVUI
Ab836V3MhMy0tgpOPeTPCeV3+TiUuAos0joIpT05W3QtqxioCXeOT669H0Uu90IDKsrNcjGwslQj
OaXYdiCvsX+5vEURJ8E6+cf0PGM5ToVTrdiqlS8MLshRwcmwaNyjzkF35cj/fWj7NZzAYHNJTR/V
yDhp9+DjhiTL2r6+3exo9pSdBHIlSzHD/NCtpNDcWd0nn3NR1dDq7PwMDF73p4wopBBNTZkA5RAi
mh8+M8pEKPJgTMrXisoS0IW22EsG7yBXgAu5xZ2tcXAhGi/ncDFK22J9anjiBtZqIfVNczTqtQnP
c1bpnfwJGeMvbhZMXPzSneIE39Q/nLXbiKg6X8DgGTqtiBkNxDOCAFM0j6bCPId8CCjkhbNZj5AS
sCzu8rpVNyE742it6sxTo+GQYJkwB4JdL3aMjh7JRCUjeCHEako8ifkO1pSUzzRQCTnpm/5lvC3y
fb1S7bG5gagiqVF5XaySKu3yvzMv8GCzh3OlhSG9gJMVRZEI3mM467kjqopKd2z8oOOMHcn/gxt6
miZ5ZAM0kcdzA/XjzDjrWDMGHu18MDYcDwRh4fd/FN3TICamfFSoyzlqzHGXJCw3H2swR2j8FyJ3
QIO3/s5y0PhqIkX/gwotXUOzXtHVcLsz4aHRk2ZluqcRaS1aiW1ndyoADUrqW4iUEkjXzzyAkfWH
GeAMD8gyK2ivIgTZmEbxh7+vl6QGWrCxqi0UwYFPjj0uO5gK4RAD1EX7q0qB5/62g9psyafTxGrQ
niOq0GsE5mh2qnPBhugfJ8q/NSnoRfmubIzhmfUe9Bb0xrVCS+B4PE8DiAuGAHcAjJQmrU04e+RZ
9JrHHzzamjAispOljngjkie9HwNNtdiuCz9Ytka71bnrQhm7QV/LHb1b6z6Stk45omMYmi8YgzrV
ueulsx9tLmZ0wLtW/FgK0nQWmZSETuGLzqeAOmwKFRZFze97apG7FQlOPHkDtUX+RoxEPOF8Jyel
Y4PXSjW3llefDTTG0ohNI8uUHPeORAKRD3UtTmUa8eh16qN7hdtB3CP5wp3fDoZz+tNQPJmsygju
C4giFuirBcdHarO5Gg6nnMNYqp6HZ+TzewR4/u0w0SWS7zGbVzvQkhlzOAdRRfxJGBl0EfEe2kg9
fSCQ3aAoHmz+1RVEYD1dYVbluvvLnvMjVAU0NBulzFkIOrtzQHV7EkTPkkhVQoci8rMApU6VIBHt
UCaO6egH5y36lwJkQXTJB34Ro6dzFUZ0fZja8pEvEw1Gtyi/PvVXvna0SJTlkKVbXZ0e2d44HwiL
ZxFCIY4RWNQRz7j5IBgb1WSA3WNXeBcAMz8esRWsrFFOZYV6tHUX0YOztTwt1vgN/FRz+1CEqzQ6
PDoLeShfYwP+DXt3DS4ofFnhXbufoyoS62Oote5ZFlTUry4R1uEwCo2WSkagisk1bMDeKMRq8c8a
hp4/eEIoPfRItSPXlMVT2tewbjFFPYPPIEzmWWHKj384XfR4Hs1rFtp9C+BJ2/1cpt6DmsvjNWw+
ng8B2QPMkqHTV36d+smRI6pB0h8tKAOPFWpOr/7ZOjclt97ejp7W9Agh9P5pde3T6Tx97umb/MEO
Ei9PmrLQ+dqtVRuJbeHYuTt7BwAgfcZ6NUk+dKRE7TeqhnFsR+b1gRHNf3v7lo5UcL9EmcvWdgWJ
6Jidr3eTXCsvqTYY/AuM8cQZtxcth/fAX0hAwRcuVMOdjUGNybGtxNjQaYdUp9KeEGwwKU3ThAIB
IxhhCNNJHMmSiEAxqccd5uRFBedyR0PB+vgjqcj9Thwt7s134lFGfEm9ZxubH4cvwk3BJ1M0qyec
U/gMCdFr420wDXtcW1DsZayo09xG5p9jpduXJq4qF1h7pINdhdeA6WUaGEy1ob98pHqi8I0JhHd1
aRE/8Duu2xCI4Z7YZFZvUNKxaDslc0EflFxFsx4GUWbMYCCgf/Ilrxj/e308Iyf0kIlgHQ4rvU3A
ViQisYYVRl59HlyI63n2WrkDJjnRsYulYrZKr6pBRDY72sqzuRHkay9PamDGBFP8zSnJDDhVdP3a
oohsGhuahrX/1nzKcN78dLRMNHhytM8DqcZxSeAwAMjNNKZ8RUJTr/BlPncUQ1iNufX0v6mYlaaS
lWhf1fJsDXjadJZFZ2Q2i9nIvEJ95b/XY8PWCw7fwOmaZ7Ptl5lxgxC9C4K2VU86SwakHJebdXxd
ij349rnRQJJ14HafYi7Pdm9lYCwCyy4Mf+HQIdSGVCNdCtKnIsT1ONJ+fsWxt/HdIxe/qoaBRgHp
feULwBMyhUGlCJKsEcGHfcsGJV78QZ+MnpAYOBHvvkQ3r/eP077/ReO5D/OLOW2h7qh3yvQ97wKY
M8liE9J5W2rJO6eThlGBs/Yi4ZOuCVCtYhizml4Vm3EjTns9acU47ODmWwDxLcDQ6+u4QlfmN+QT
V1KKn1ncmNTb1OmrxBm6Xu8Owgc+9CehNppE4RT7raDb+ihsCRO6MnTiq741Gnf69D4oGkFq2eyb
I3cB/d5H6eEDxp9BxQqwmqL9NkarHNU+96ykFP9DFaVDm7R+2nI3Pmv2fmDIACXXaRCfiPm3RRyA
iXYQ9ofDdCky2a4cGkRam06u+61+WhZgu/hXo5vDY2xHC/MSBw3mX1rwsGCcBEa76VEk2TWkJjzp
0H60YQ0i/QjgYkwVGGj+79IF9y/XPwQ8HutQI74kk2xZy3kwxwY2jTkxurRGu2jXPNvJ66QNhG07
kCC1M9HGpSpecXFwkd3TF3x919JXPjKF/+ABl1mC9Yd+EJbAugIazAitjazLFJP6QVRQ7uRlHIiR
KkQFSYoNy5b9RQmWlXgrUsU6DqUR1uDPEEPnl+R+oFuvQeDcD+1XdXiq9cRPbC2DDvFjGTe4wG7i
bNMJfX/ZAz4JudLZnRvfcwmSn82h0e1IleJvJxLRh1sM0FMNi/zrEiMYYwzqatl3MYWn4vM02T6n
Ednh1dAftehgDU66wlFZbvUw96PWrAu/o2N07AcsEQXqrJF3LXBGmRoxd9L2BcfOWHWVfOYn7lkr
EJQRDgkAOiMma6CXz1esfD+y+v3/zNtQN3BGRVEP6l1uYTyID7ZCKNd+Ux1GD4/cuBdhxApZmeeM
0HgUwFpdtISNXnTSdT3II7uzJnPu4d78vyT/aPmli2TANbt6yMJBIcXceWVlRCN04wehXfJGqsld
LXSV/pMdMII2Yk/ZVP/ayGHZ2l+LkySQBp43pCkvTRgUe27ePAiijktSvE6YxQJGHinw7wtMZ4Lb
eO4KUfjMHJPpgc191Pgh3PxAEaPSOqa98vsTHVCf9CgdJTmr1hE4nKBGXzfjef7Um9XaasQ1KmlD
KfuJ2vP6Xs+AwgUmDN5zSEdR6wuDflHYHJ4DAgIpHT2KNeHMRUxtQV9Xd398myhl7+TwFSIKP4/0
PXN/TVCzdqGDgiRgGdyArXK8m6BVZSUkzvquHsXGJYtONu80vtBOnMQs7FKZq3OO2+gzBwnfDdMM
yiuslqn2iOboEl5uspnRn51BUfg8maLdBnfuH+CnWz8+kf0tRxHFyQZI0zhD+SBbiYxjE/eqt4sW
UcAjoi0Nb65LIzhK0PcsVKEuIXicGqhaMEfh+vpFSpt4KJ/gyJlFIX2vGtC8J/EpkOUaYVIVilP9
RhM3Lm7B7xaaZA8h3KQR8wyjm7eDKbW0IxZnFntoOftNib+oSDW5AHGzGv9MJf6kQ3RRcFCSb1qM
GI+0i6uwcEhzO5B3xuu78T3OAwj16Nf4PEeS/pQGJSD3X1DF783Rn32An1GgVsYAcJ/LCwXin8z9
a3/+jZaNPbbVT77TrtETJtvjNj3+sTMbtoFWoKmNCEXwBVrTbjHsmRE1e2lyJF8VlTWuqDJKCsdZ
bpd8yxDoyvClPkQf6KzJF60TPxWiGCCCtSxoY9BPmDpNeY4FUyU0KO3+S1mYxPim/l6N9WJdQ8j+
O1f3N4dzat/U4fI5Og/jRiJGD7Dn3C7bGKT7za05sVX4X36zdpgT+y8js1bz+DsdRs/TeIcs0Cqv
c4F6KnC5hA6YPzBLWd1yqY8cpvoxjjuYc/JmvAn+Vn2M+b7u4Y88euHyouJ1p7jZF+UPt8yLVn1a
ozie9Fzjvli3SakZDwsRxW9gXgoyzu6VwDdAME8x5Uq/u0vsr1TJERE1N5wS4VwLu7YvMCBt9q/w
ihVpu+TxzBr+igIaG8TJWhvdrzgWnYMKkpXyqJiqz16k1ffAcgWdoP/ySEF0P7n7L624hubXcjtG
cjZRPNC1bCUaRcD824yIa92kAOex3KAABmkdLrF3OTic7hmnF4sY5hkPM0+9xUSdH161BVx1simI
ljaPYHh8BT7n4XzeT3bzvlczcVnxeDnf1mSAXVMfdo8tlno6EZV9orLVtsCVIdi2zyeV/0qF6OCj
FLe6L8aDx4MQ6jAWo2/eQVQ+uh083Zq94gZMAYrPW9vKlbxxqSv+BpNYj4DJXMYvSA/xjVoHE4Ak
JfBAp5wyAckHDu9jdebV4tW342bvrnQqW0EJloIGRBsgsRM+5Qtpk/8FhxbhCBK3kRyp/O0x2aCk
2fZO0FZ/1pK+/76Z7LxJj8m00eSjdliW/Q1+461bUmXSdq0uloQuwVHdPTXgiL9QNKPU4vlDtcJ2
uACZ2Ou7xiNLEItV5IwcZeRkg7MNRCC3raTmUMhyY6lueGmvQg4hv8lv9dk0cNOSMk3f/E9UmF/J
j11WZIDCD9me08OTUStcG6a9FyJMjeWgjqOiO0uoAWUjknNG5Tz//sx2NTR7ctHmGuAbG6yyazei
DhbY4R6toSjuLMJnpXHgR6j7irxzwEZWSr4HY66GLuoWr1oTK5DdoLRwYbXyHFN2FzZ4GyYXJXGJ
R79bRJaH39Q9sLxiz1WG82lps/zMMxeHGLmCbtpPusqUvSHfeGVhe6nYSC4EOWLfNPg29sPRi3+H
lRc3J47jd6iWv+P4qo50JriNbQFnkuqWVsy8sMoIEQtugwz+7AihejeXUK1vRUGDFm8JYDLfnzWE
cuyYeRCT8XsJu3YmuZ308VJMraBEAkMdNamt+EoPlWG3pKxWOTYaYg3CnxSAoErtujF/pnMXRFTN
E0AtLWzdmfZ8SDqvEVRlcgu43VY8GJtkAlz9CUvo4JkigoL6NDAwRUgBwZ00/REynn4VeuVOEMPI
HWjjQRNQR34/AYT0xnOmL+pLjhYcJouge45oNZ8nJc6kvQI1IVvpJf37QnEpUpteIzZM1b/7Cb99
zZURLEC7H52tSgsJQ1BcEknhgBhy+8qeKQxlfu1nht9dao/GC0r1oKleqxviBZf8k0o8uuFflNkv
+Ue3zQCbPz7zMlvtVZsYGaj+HUYcYppQRVVwruqkXrypGsAC6xsaJBq/wjsWRAtSm6BweuvrrMTL
zInMYwn9I9nwZAWbiPM3TnW+raFBhkbyhPzR8b0rvKfOlSOdastF4vSdBwHyIdZUM4Rzi1o7KALz
pEhcjhrS6bn1RrO4mqQNs4FwCv5G1wP164whoW82zAX3li+bmEBSpeR5W3Nm37hBghIVRZYSLOJ1
H8fK+DhVVnI2v439LQV6qi9mGLnQGudv1qyZJliRJTKHPtlr0cz5jf/54twL0gzycS6mEWvzjoeU
HX2ZCisbsVyQahvHgauj9kM5uzc0yJlw+vl0jcl/jhnXc+yHZFyOsM43mIgufqWjQo7k1G6VHRAS
uQ6vcy8Aw2bmOi972kF9cq4VrZN3d7HrAMF0wTzwrEOxNKR6KZNPGak9YDgEvVt2QOBw+NoXJ/HS
Ud2MZVB/+G2AcNuqFzff2J3beMHosB190Fqtf9z12jSIbY2EUGUqRdSINQ4/7gxLiRU+OEHpV8v3
gOSKbXpDOJMPeOq0jaVvsxytcRjuISVy51mJ7IqCtESutd9sUxxlXtUkCkWLuwl9WrwtwRUgNhya
CwJaHXArmZKiMAnpn9A83eR6Oka46v7xoxnyuhCRnZNpJDkMgFBxiaTK8BDYlGhjnjaaxlS/vUhF
jQAvwbgEDvfMka0jWu8Zh3246lTasVh9WkIikGgO+jjgFLXngiH17Z/fM3Q3PuzkGJxpXAs+E+eY
msERuj8onGRe06s+r+/1o/PuSgFZy0B2EZkmkWUlaQmlAq3hPvpREo4vzV1VT+p0IuiOe87pv3sw
jiH7vAB4zAMN89YuoANY2/ldY0ssR48F7GEpn+ef3jW8BbHY+ke4Cr/Q8zqgo/DZZYaC9Uy5dh+k
otZ9Ai4sQIpJCxJXLmV1kv4EwmzdP148AVKtuOADkqWu0RjTtYyLQDLVC4yyLhL/xr9E2HYjoh6w
WTyPmnrKDnD6h/NynJdrF6QP3Tmx4O2iE5RZSA7/3KjXWrwfwJ9wVp2loY0f5uLbtePjSLSBMeHg
gtIVuCCAzdDWNekXPce5dP8nu1R4NDQbJJBm8gjir84P09u/jdo68jzAe4QJkB+BtNPkpRqIOnha
EzuiVdRPN79zYiFltSOliPVf0rDthZc+Ji70FIQkaD2nIu+pMKWV22LhljRR/bkKilkyQ2RZlEQ9
gMk5FDo6n14fFf+5mhzic82XK5t2tpkubCFdcLGqiS1Ecr6FQ3Xj8+pd/BWWbngTePGYsLHO3T18
PWfvIRRNaWlEZNNaURe9+3IX1TkkhtKqbHg7H8L3Rnptnht6DN40YLX5QlbPikFT66fVgR/Nuap4
ONQSinhzqvPZeHcwaE16ZflL0qjoljFT7l+OX2HgpBXdO/T9Ibgh4c65prsBCtTqwSdQPXlv5rUW
j493fMrv/GQgSag0YnkJj/JF1dPgsFznzY90YjS4a3iIgWC+8k6KbS36zx0i15FVnjiBFTlNmwmG
9R7pDuRLfGXAe2OHen7QQ7awxnYUCMlCaWU8x/ucdsN3L2odE7urkYK9WxUyRoGIUcbpJhMdFDiv
19uvoKdIOvVGL3q/7cnrbU+Q8eaEkycZlI5NG8iZBiBZ9m84V7ybeOZCxcduhujSeJ18rRiarTlA
K7ooVn8uyJvoes9kN5aVP9SxO3Hl/bPRIsHErGdAVw8RpAtH14jw8WfZyfTmsHigFksW2Kgqo3hD
eEl9NP2TsHT1L2jWmqyaOXOgZV13lXMYTKom+s98Py2aJYmmy/KFdMwi1/xxNytARv3ioz5UEXUI
OL19dP0OIKThKt8Jp6kvdXwi7wtDbLaG9YbB6HEcYxroWEE1UGv63UtjgtCuHFPQ6FpFkiHG6H3X
+agcrbnnLCUXR1u1qDMq3RNxTIuG/nVGS1dxOqNLfSvafmhg3inqha7SIaG9erLwrov/QDB2VRSy
xKxit72oWDgN5rHnWuPiOR2lHNMcBfAgjvtjOMuT+9eEG5Ff8yT4DqJVOF1go6aycpjfWvUdfcKU
sLDFl/iFN3RlpI00WH3pZLLW9rcwcNBEw7w/l6sjfcb/Kts27lNm1LiOfGzUy8cGa/kJn3CR4KDC
QVvl6DGDBnpIEqT9P9ukChHvubs4FYuS9UKCzdcXDIRdldOBWf9zse/Ree7s/ugN/ESJbhQKqAsB
eC/bn/EYmJ8iMoO4wEi9KDmnZ2lb+Xz2WbIcUOp17SoxjCCG4NnLJ9uTZV6zAaReCIwIWpxuU7Pj
NmHhOtpYDRSBi3f/lZjof5zSlO5eSD95uxVe+tMeGMaXdcCvElAU2xfc4L/2I16sZL5RvB4kOnQz
Di6yG4igg+YkC3Sw4tQEAfhpEOaa6ZtmFTDndju6SyowEBIQ8roYdsUNipG1nS7/kdlvrgBV8C4u
aShb537JgqpKO5oT09RkUk/w/Sf0a/D0Q/FHlVzuqh+W1D619yt30sHFGtFOTzYHsoFMaCcrFazb
FygRqdPrQf9ZI0ZQMZG6vAtgJYQ4Qd/b0dMdVmFMgXDAr4aPTemGMg+80SbtoPUNJ3isvOxjYAMf
Q4UgMcrxbNoBqmVrCZqcgPKydP19o8smQXD+8c4MYzyeBxB7EcmMmqTRfTX55l8RsoA0+eF+sFuk
LZ3efw9gfvJwx6TVOyZv0vYF3AC4IQEcA6kJnZsFWBXzAf0TCa/sjtv1hLX5GhfYzQsAuhZHs6fD
sIFZmcuqvZuxkGaafwBMeGsTnQHaA4/Ncmjqz7NNt5qWX4osxN/lW+OGEqM5kZb3krLN/4yalXQI
xk2NmezNZhWLxSIfm7zVGgaWtRhsTnkzCB1qqJoLeeGfuTC4XgsqAhlwk7FNR4u5USfymoz11GtF
CfsLZk4Mr6YZUFFbsZzouhtCMrpnUM5ideDJSL1RUVS839PcoNrDPVEOJ5q94BqgGmL6gL93noDp
7nKQ4+kxmmb8Kl6YKtlNEWyFIZ7nXEMCeLNdQ166g+Xc91U5QURbBglHknBbHvnGkMY5GOlbmNzP
/u3vi9ACikAnEK4Rj3WqY34/1imYsJcgJU208c0m3Jbihwj20GNDToDywOskOygBuWMsW808GVuO
/F8NrZ8shPGqf7qAG9T1TIdvS/zoPPgY25NPkZeEvnaYQUr1edyh0/o/pJIpz2x07R972ZyPOTej
BB+/1R/du76nl2iqud5DZVnHcdauxnFI8RWtqy4Cptqe57jpWLDE7HqLO0U4S2Kj1r+tzmj+6Iot
HmY8WvzlabdKUb9F0yueJ0Fab3UwzgKNnL37rNXj+AxRFvZS9nBDmMGtrsEGOyh+ptrpccQoswNo
+BL9TQoGooNnWBDQntCe648Le5tOJsVUHSaRXzzn9cgErPHxPaaY8F7xAfwxw00JRGkpo5Manfwd
TojKX6b1hbuDiNfOPH9j5fp9AiT7DjFo1XxRaoZZ9oHuzjSzZkva11xALAZFPf90/7nwp+JFvGTH
EpHb/6hzGFgyLMZ78Lq8U5tjeBgki3YV9Hoy+kxJsmNKsRjTLO9oqetBQ0VNzvVYu+P/k1iGRzIk
B6GjGDewKtK9y8QFF1VS5lajksV151UdA0tGWR1x4+k1EWrX4h3xgh44+3g1iToTOJy1NjmIEdiD
FgCd/JeRQmyI0kLBPGhgyTj+SNt7aBKB9vKx81UZILL981HNrEaJZnu5EGeeUDQa4jqiYm//WmWP
l6Pa9yzxrLMFCHFbUzIJgmROaJ2809iLrxrmEKY/Cv+YbVqs37msWm5T/BoNtue3RnkjYCQHWjxo
Q1QX7vaviaL7fZ8Nrt9s6KLS+PCvASOZqf9iXQbndmgXyJdk275pSZyt5sfEZ2s4TQEqoZ03ZX24
31eM5pLOReCcfWTbg+vT6NO4fasnnvpeoH4JI+o4CTIiWAT/0hUFARJacJ4=
`protect end_protected
