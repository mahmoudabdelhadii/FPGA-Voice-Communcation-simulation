��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��,�y�}�ǰ�=4d�H���`I"��W�`r���T:tB�T4D�m�)�	1��I�t��
��8(�8t>s)ו�."[�漆���]�~�]��;�O(1#5���D���d3�q	��9/�I�w`W?ދ�S"K7��5�,l��C���
@E=D��!
����荾Z�V�h��c,Dt��&�����]4w9K_9O�=l�uE�w����[R�\�zÚ�-J�$����åCj�[�
����T=���K���h�����,������#�z~��?�G���B�~֨1)��k��yq�$/ju�YA9��SX�{@��mWt������w�F��r���������O)�mC�&�����$��^_��|�����=������A���_"�s���50��-�ݡ��kVE~�cu��'Ah%�����v2ݲK:|�g���7/��=Q�u�~��qC���
qSa�a�n�m(�]�h-�FK�]�Z<��K�b�s��'�����C$Yכֿ��h|�[@lXJ�*Qm?�аR��(�v�vlr�j)ڦ��0p�s�bv��jy�-����(��N�vהS��Y�n)!��\|9��;#�o:�#��9|TWL��L2=�'���$ƫ���19�?�:H�A���T秧���,rJ$�p}�a�ڡ�rn#9���~�1e�[e���!������{�T�7���O�z�������쉎�<o�j��D�7��lS�ƃ���F�V�:¦?�,�:4I~P�o6����2
�ԫ�#��G롔�qH���'> x������>I�nN1.�yφ�V�ǹW�)��	�3���k��c�Rw�buRA�8����\��L+p�����U�|4�}��3w���n��B�2�Y��Bر�An;|ܿM�MT�[�=��Kv^��L�`.���kS� z@���Y�'j����@ڑ�Z��1\֜;���z{�ړO_�C��m��UW�˯�1\���-�P�DE��`���_Z��6��c���꺣���ĩ��~ר�-�L6�ɜ|�S[�/h ⲕhQ3 ��Ś��u�
�6���;�+��^�Ly9L2��B+^��)�f-µAE�&��o�C�'�� X�a�Ag�4����R��X��@�;�D}���|�"$�ו4J��kˑs9|�p�*������kIYm?��.=����S��2"�Ѝ�����/�9���M�s�?��>�?=�7��V���hV�Ws%q�����i&`�B��?81�.���󇏊�� �#5�7�Z�o��r��no<b�z�N^rt���E櫗�|KS3�M3�@��E}���6z�t���!�?�m�}����렿>{�{�W��B��>���m��nm������ �x�<1`�6���G�G�w`��(wΖ�U��$�ju�AQMJ�4 Y�d���`��h�0�vvu���J�23(�;-?t2H�y<ǽ�vڴG�Ji:9��<s�� R���h�|��4���E���z��I��F�@�jKFB�g�`�}q\Bb� ��A���n��l	�կ��'���z&L�Fb��8
�%�a��|J�@�l#&H�
��o�
�3F5@�C�])���Wz��S`���/ ��?�rAg���B�4y��_WWb�'��8ֶ�<�ع[?HE^Ѥ/�ZJ#h��8r9�A%�o��W3h^�����˾��Q�;k
�?�!���A�I�c*~𴤊U3�ٸ#�����s=��`��<2���1�t�� ��)	�quׁ`�����]ml�����3\l^�˒&cD��eT�r��<�J�>��*�~�#^Bk��b5�7rN/n�V%pi�C���(�7�] X���K�C�B�h�� �����Hʮ��Y-Jaq���QZ�(.�b��Bg�cSm=M�ER��T�ntB�@oV!��U��
Y�s��%� .`�7l���5h	��,�#�%xq�P���Ż���f���IX�:9�o�ߝq�ËV]�2b:=$@9;�<��\�8yP�(�����x��Q;m�S2��j��j�P����@W
U�90҅��Q3�d?����*�pX\1k�0B}�;�C�k)��4>��'����o��U��o�Vo�V]n��i��^�TqpO$3��+#l�4�Y��D#&�*47v����O=/b��+χ��0
�X��V�����c����ܽ�n лb��{���OP�	��DXDk�G>������R����uؘ\;�q�ݐ�8������`%�P�x!Ym��#b�'���,}p�k����]��L��¦���\mmu%1,��,Iߡ4dٔbn�ѯ�魫v^�.T�7Н`��)-��p4�.X�?�����]�&����� ���F��]�Y�>?tb8s~�s���2IYe�mQ�GA�V"g�����n��H(k(O+񸟈�2)�N��n�d��k��C"�Sz&P��ݹ�J��\�b�
�� ��/�"�D?��2�g������{ۿ\�W�ɰ����@�6�^�Qz��a� ���h�V�\�1&��T�f0��ia'�S����~yvQ�RXJ�F���X����Hr$C��Z��v����mb���]7�3�&&~`畾�w��o�
'|G�p�<O�ߪ�+Z��&Y����v�w�1�n�<0�a*�瑢lX�Up�9�}�r�}��]���צBu�m�2��ˬA�K�` �Q<Lu�N��)R5�H�#2h���~��	���J�!|ߏ�����ɤ�_%áMď{!���i�&@�b�'�w�����s��K%��� rU_L���s��z�`��=?��𶦹Q��#.���5�PsT�t��T��4�\0��6J�Rօ�5ׄ���S�Mo?�����L����]����%D�(C�\�ku��|��f��!m��.܊�-�Z��m3p�kn�WH����Q��a��i� ��:]4�YD��[�ӖE�n�{�������ˏ�zpI��=���֊W�A0_���Ћ��>o`b:�&;EEu�(L�Hȡ�k�vŢ^UA�|�,�mj��D��1p�3�E	f�>$5�.J�)��{��Y��%�nd�����4�u�&��8��4B5rNֹ�yHj���v�ħ:��y�K�4�b�a�oE�ed��A��e]64����`]p��4�o�ᵺ����B���Eq��j:��:�8�Z;��9�7w;��Jiތ���E/��B�8MH��w�p%G�V�ܫk���61�_�� �����v�+tmiT�>ԁSC(�@T)Qͼ�b4���$�V<E��\�:���2Cn
�"m�(G�0T,0t��O 1}�NC��>oL�$�K�
	xǥ�,��&).�g=�tV�l�	��~�m�y�z#�e&�wПÙu\�D�>̲:�g��Z ���#��
���@C+��EVBԬ0�`(��L��@7����_@͚���'�Ͱ�/�,~�=�ݔ*؄! c���_�De��Ny���Z<YC�o9!"�����8Ի��EB��L�#� I:6���kt�Uk������A-��j ���f)�sⶴc�~04kK�cL�U���L���~���*â��<�$�SJ����ٳ)R#/qѡ_����1���Qt�?���7RV^���+n"b�r$�@4�+��@t�a܋@o���w�p�0�ş�@��.�{-_ǌ�����U�n.76�Y�	#��}�t�!Z���v<��j�85��IŔW�PiK
��$j~<���H�0{��0��L������:���$�J� �ύ�Ta4, �GRN�A�sB�%�į����)F�
�