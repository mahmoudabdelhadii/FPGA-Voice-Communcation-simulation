-- (C) 2001-2016 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
obt0vWRvd/Wd9sUWZ1x8iy579fGx2ok1PrBGowFzCypSHP6CmLS2eH0M2CVJbRaQorrytU1C8pFP
yAdllEdX+rIiVP0htndH6Omf+P8xfjTVR1S3dcJXzqWiJsZArO41gluXxGh65GSAeJ+vCzaFYsXj
zcPT55v3ffuGdBHUIJMj5EGZfi1OwVe1uNYpdI68myQ4JXf0H9tl4RS/t5wyX4QP2HXdq0axm1vY
5Jh06pBaJn7k2Avw8eUMfZKaqfBWe16MDvuEtvf4LDuhrLPOlaInAWEMDLXzHPlpjNLTtvamlnEp
vVYSMh+XB/P3WdH2y4kp2qnN9+yaVvgyGMn8Zw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 3984)
`protect data_block
LU8FjKl1qJkZK/lTlKO1MvgNJU9KFVPg1nZy/UWcnYbjYsatiyqLpebaeDfEKrXYcre7JJOb/+Hk
bIZJyegAmyhj+mVAPeePC5SKo7MI4ULZewvrwhmaViA3HyXvruYlktfrSssZ1tMk5kFlTPy/3v+A
Bw72brgysLdgjzo5f8VfLo21C1QNcnBz+Kp/J4yy3/aq7XwlB7IZEDQVL0cYmMwp2LSTdFDuhufD
W9xe2kICfGLyFu27WSfkCSJfdCfNnTLuvr9k/Nn5s3A2bJRgg1pOslLMfi9DxpKZup7GQdUHJ6hT
+MlpACdTw8nP6OsnIz8G/v+bY6CEq3b+rcgpM/pO1Xuk/1T7K0UD1kypz6FhbnNEYzwEIcE6OsE4
7IeBPndARzIdm6CsPh079aIz7WOEt1ak6w+T6+nP/p8rezJK/TuFEMPweKe/kGFSFIsBDnDjtxad
35YMxIRXYuZ39oDCrtvO8kGQnT2cGh2DR5scvxKtZArwAsvBNAx3USVlrovFzqVDkeu9Y9kJBb7h
h4NGj7RPHW+pksnHKSb+NCn6un0FOTL67321ahB/6lGJ63c5Nq6yaRAr4plxUH67ya8kyN2cbe38
y5PVSTIrvkd8I1fyvi8+EsWYFx4lt1327nmBhfmoKp42IbleE8eJ1EqXaToRcY717A1hqMBnqrOf
5hujHQ9ogckDzRpc433L52Ji5+XWgfVCrq1i2/vAI4O8FOEA5OxTaLbk+VkXCvZUzuEsN/akAmiE
BJ6cHzvLKzAxSgBTvwSOBIxNQxpr1wchHp2VfXY7dKEVwSrpyHBUmQ0w9zIf6i6lKR+ogfCAamB4
miB8XJB7sGaOsxvcvgNgeG+F3WNGhiJ6AXYFcbj4F6HO7fMzBaNnSCyJnLm9kOYsU51O7lcslOKq
s8NVraTMC1RjNRe4OG7siJGmN9a0jlXza3YQzLai1Vd5hQsoPVB3THwk+dD3Ykix+vrvwy2OaMyA
Aq6UBaHLJsFvPCzZEU6ZukxLtgV5jeS/xdGzSMH3y21/WLxQ8qKccHP6BguzlSUe6XahN2mmDc2W
nB44tAl9FhsYyuhTdU9HX0fRKvw3jY5YfKlW69/ebLAlTtIGMckczuQllqI96dhwnqx293sYFiVU
TEnK//WLxi0ClIObyMUSd/b+jaVi0dASqldIq/FQkXLeVOxq9hloPsEhSb50AcVPm1dKKcMZT1xT
4ziVAqCGm5ldTB5lzGGNEeffvC9cNCXgFIBZxl6OBlf6EaO3FjCLqZWYPuBLxxm11w0U18KeQjX2
YDGpdBQ1v82jz+fl+WgUKK4BS8i6evNv/WI42/aARK/fpZVX5ZgCmqOIxTB+LdoTNisjq4htzCxU
1oj20d//+1TGta9+QMJLSFRGyKlZ73VPyctaRQnvFRQo2J6B7BO698yud+JHJ84ISZNnMl5M4/3A
kTQkwyWLDssQvxHlWFirUsiiJtpXGTFc3u49Z8QWcyNXNDpY5I+UU1NjWQwT67FThkXGFvuqgn2E
EcHaFipdp5OHrmCDcAaMTkpuZJoeRRFSGqg3+h+bppyPmqQUNtDChyY2+ug9OIqF6LvZAjd5QCbe
NAoRh6p5DlCxPqhZ8XkC9s0FH6H7bTaRQ6om0mrDIjkb612/Vh8q0ZhpSn7mUw+z8K8Bjobt6MzW
xlC3VlwSAD1rRvTYEqa8XkVQx7Tl0Q5jO5wWf0OhtIXuj6OIhQJEoFN7zw8wk8RTpRWmWouZDUyG
zwXqDJBoVjmi0rTePyOrNMmKOnnvQuS6WHyM16TewRNbOL8xVpqY6xU6FbIJpFOK7F5cwxABHHdS
BQDTPi3gbdMzK12eJBpMFT/NTBPXsd+y3M89KxDbhLN3ANpNXwwDk0uOGuyA6hlvuRk6+3wWDxe9
7Pb+Rt0YYU+G08ykkwfM8EUzqLfQ67xm7JBOboyFrJOg3rEwbgW1v7mEqDDPxoOiostKIgfDg4fO
Or4pv3gudWkdes2xFCsc0gyxmhPvwwmGsFSZVeIX4T6XunbAGLOdBd6bCZvnbxrdmFwlYwgiGxSQ
ZI2aUIO9hz2UFUZCI6SpvTKpRT9a2Ni0u1If5aEn210UaXetZFLsLt/20w3mw1N+Y4gcJyxHsDlx
Nj01/QkfyoDhxrWYFWFrvs8vVZcZq/NOMEswSFnnvoaGCl1m6mTYqcBHKODcXQTmkEpK5p1D0dWn
5ijgyPELNhz92ZaDHcMNon0aysnx6QEPHoW5th/K9baGb2D8zbTjYffCrdkNfab+TcTaw4ebJa6i
F9AA70emibKbo25ITfYRK670D8GDvld/WwAdJ0M24lEfnCEiQ6yx6F2ClS6A6gnhLXheBZ2QwMjd
6wDliJ8pSuPmPL4I9WNsjovfx/fCj0XNe+VqSDm0Ku2GdKRr6xnQL+INP57mteeIFtXPwXn19u4F
GQaBvl9JYPlrZGX3f3QbVi8ihp+uEo3RN9mQEBpjEr+3vWkdLAxLZqQm9MjuWOLdvZBmXztbz1dG
NZlaHnWy1YZOAPjYzvxpAX7s1Apee14wW30cHFghsIgdnYLtS+RX4w2s+W3b7VmOO8KtUVAOEWyi
UxrScA4eLs+eg9bp9feDAXUZiHn7A3xmoZQepnULTA7OCwTuXZKNlPmtXQ8kwEafsZaE4tMRiiZE
bZbV4sQxDjMpCAEobSKuT+6JjqMZWz0U9AVLbAqFoxF9CYMIxlbzYJeRyGQdPyncEBCS0EuJN1xu
zEF1uyrLRHaGG261PDEAZOJdznVeVtHHpM86dmb8zkTGGRm/E4D2BIX65g4T1cw2prylz84oR8iv
ZDHHyIB76NYHROOD7KJLHW1FZvngIhQAGJuYOseJ24SY0Yui732A4t8lG56eFc97ip/wdzxIHcL4
SEaNXijyYssbWVLeI5JxfltCwatn/3Y5fyNCQ44wQL2OP2RsRaEsUqBs6oO309nR9ewFDFmHrd1L
8pjTdwKKESMDkj/bfyZDQamvxcxj95DsHTndpyAEUBT2yOXV+9xa4EZqM4xJb55X43mp7hmwDx3C
XrgVsEsf3V341Z+Be/zIQVhYwMOi5yv9WKrBBvTzh7cqPS0vGpU30dDzR6XQqHywYbIUsSC0VCRO
cS8NUxsNVeNzYdXrFlgI3lOTZ8sInfbVhQBK0ckClIhPVHn7Z0rG0obL3fInJOm3ah2lEaBBA/P0
XvKpjfXb/uFtuiKKeBlE3kPrLfdpXUR3y8v3a/+6hnZlzeuSLeYH3//+rQlN/PX1iRA6Uxh4ljHz
QgsiSX5FqA8YMXQ4rnrOnbeQyMZ3kp4O4afx6cXlWTMIj2seog1Cj87wutVqLmTgJMNkZcBvzS+V
xutu8CCL8mrUCIuiS47zcaXuIXj8LNtME05KwqZe5sCVsU9A6VgPlnt5blaZR77Y3PzUcaRngucI
/+gRPPBu4SlocXIxz/eaOlaa+8bjJnEdxYBq6Yl4jrvl4mqw52UmWFCMSgNf3ztEsZTFjZnkBq8c
7A+kfb8tJsfid0xs6J3RUV7xNaf7EU26b1CnTaACavqPDG693lrT4a8gw+jBTHDs9tLAmvH2tL4b
1h7xzbQUtgbkUpl3qC1b8883RVr1yxVKXjC6LHrcNvko9x2ykb4r22wqNLwieLgKIX5fxlXcbBWF
BI4cd3+3/djgBMDFghGQpcufKGQqCQY5Kcvwpt1LKWhoFytljnxRzxI2XowkDzN8qHsLjnoa2GpE
5cvSIiE2TuhsGMeBSihjSbPKvOjZ4FAWvHocQ8ijmirKOe/xFyi+WWnu+g+HSdOTeelg+HKHOrym
cKIaZn1BfSfAaXupGUqb9M8g+pci5Pwwf1PB+6svEWvDSwLqEsznPnybqzN0IqL7aLiRD7Yzzs03
9uxwSOtOipcFR8dRetO70t6ArRcgCWlypu4Lw0m982Ia8pSw7fYnQnQsHcXHKbJtf40NZXWmdki4
qqpldN0JFL4dgR/whrsaoGfYbF9D81RPhy8UTnEaZrKeJV7ylz9j+d8Zg3O+VejK7o7X/u9e+kkn
wXkZ/Tk0vtoGTsWpDcyziLhUWU9OyyeEZmLrPGE5SNovmAEQGW6MIAop65wuPt23ZiC+T6nbDSV1
TshGJcotj/4HFwh3gyNqjGXCrhhDdi3wZ9Y6bAHKz8rayHBPe99MU5rasRVeJJBT2OOuxFXHVotQ
ffaur/mK27oDG/iR93tN8s/4jUwGLThGH2I5AsIldIqftNFInw8b+OFqCbtI8Hwzkpdc4VUSwjKU
0as+mp8bl+EAzvcgiJC0Vrs0KEUi+OQ+RpMbgxbFvrfUlZaeznmDEDwMjeXiXNZ/+Zr/exmGVLb0
igXTollLN6zLjNzISENx7Cs3dn/BYZeuxDipGaBzwR4ti6v/pnq6H3jruob6TXoiJ8nYGCQhSr2H
bndQMO0ez5+cuX5uY33bYcGa21QjS8tHqZFihddn2Ca17rPGm/lgoQJlYLcno2Tl44+SMnLC9lZC
r+SNF6EH0gURz1AFf8YjUKpLvmb3gXVj/y3tsvZtk8EdGD/5ugnDVLhcm3XD78eXMu/oYXsxCwVP
lx/+pkMaeczOMDznNj9DuG9FqStnnHKXV01pFjoMcD9a2fG2Xg2lTb3ZrwENDL0hOsa7ED7mZlN9
sV5DZNo6isiIgrIiuV/TjCrVxu4WCKPJ0jR64J2MsFw9rW5WW9/qQUJORN7jSVz7KQl14Uv8x+8Z
6/aDf3QhDH5cLzGvkgFvc2BkZPydQXuw0JGkysAtgI1s1p099jQy98IbgfekWvyJbcrC+e7o9XET
evVY0vMrxzCloRCkny0htiyIfisxeLj9Mn3LXbL5WaBzRzwDVNIykCjqzdyiM7xYJuOx+3g0G5dH
zkUXeP5mqosAVFdU+Uy3LhAPXu1ggBZcehgUakZs41ITR70mOawz0ODbZoS/mcQGu2fBvkZl1hGI
kUEiDpnHPeacmhfNpzTQvGd/V4TW1zQ4AVhpWTxYj8RH5fxSmwJgNks7XCR8eYLQmk58C2MZXZgP
2Jb4tuAfYw0cqCncRYaQP7zn1NxVXTviF0G6579U0LT4ZREGHaBo76qGyld40l2HIxIdk8e6qJzm
CXyVNl+KKUezt3MGZnu/bO/oeX4uVZdYjJAz1i4h9ayfVCOzWUsbee9Vk4AP7P7CoP9RvC9TFynP
ErD0c2qmyhU1e9orTs2PgSt+pJ/hFkDegKAPvgeDRCBXNUN92SVvUebAcemyq5zhX6dZFPImj27i
CuTVQUYprf1E0MYMdxtdUOw4gAzo4kPVJp2wHVLmNR4CGzjovMF2tsKiyYeh5hMMTrjS
`protect end_protected
