`default_nettype none
module Final_project(

    //////////// CLOCK //////////
    CLOCK_50,

    //////////// LED //////////
    LEDR,

    //////////// KEY //////////
    KEY,

    //////////// SW //////////
    SW,

    //////////// SEG7 //////////
    HEX0,
    HEX1,
    HEX2,
    HEX3,
    HEX4,
    HEX5,

    //////////// Audio //////////
    AUD_ADCDAT,
    AUD_ADCLRCK,
    AUD_BCLK,
    AUD_DACDAT,
    AUD_DACLRCK,
    AUD_XCK,

    //////////// I2C for Audio  //////////
    FPGA_I2C_SCLK,
    FPGA_I2C_SDAT,
    
    
    //////// PS2 //////////
    PS2_CLK,
    PS2_DAT,
    
    //////// SDRAM //////////
    DRAM_ADDR,
    DRAM_BA,
    DRAM_CAS_N,
    DRAM_CKE,
    DRAM_CLK,
    DRAM_CS_N,
    DRAM_DQ,
    DRAM_LDQM,
    DRAM_UDQM,
    DRAM_RAS_N,
    DRAM_WE_N,
    
    //////// GPIO //////////
    GPIO_0,
    GPIO_1
    
);
`define zero_pad(width,signal)  {{((width)-$size(signal)){1'b0}},(signal)}
//=======================================================
//  PORT declarations
//=======================================================

//////////// CLOCK //////////
input                       CLOCK_50;

//////////// LED //////////
output           [9:0]      LEDR;

//////////// KEY //////////
input            [3:0]      KEY;

//////////// SW //////////
input            [9:0]      SW;

//////////// SEG7 //////////
output           [6:0]      HEX0;
output           [6:0]      HEX1;
output           [6:0]      HEX2;
output           [6:0]      HEX3;
output           [6:0]      HEX4;
output           [6:0]      HEX5;



//////////// Audio //////////
input                       AUD_ADCDAT;
inout                       AUD_ADCLRCK;
inout                       AUD_BCLK;
output                      AUD_DACDAT;
inout                       AUD_DACLRCK;
output                      AUD_XCK;

//////////// I2C for Audio  //////////
output                      FPGA_I2C_SCLK;
inout                       FPGA_I2C_SDAT;

//////////// PS2 //////////
inout                       PS2_CLK;
inout                       PS2_DAT;

//////////// GPIO //////////
inout           [35:0]      GPIO_0;
inout           [35:0]      GPIO_1;
                
                
//////////// SDRAM //////////
output          [12:0]      DRAM_ADDR;
output        [1:0]         DRAM_BA;
output                      DRAM_CAS_N;
output                      DRAM_CKE;
output                      DRAM_CLK;
output                      DRAM_CS_N;
inout           [15:0]      DRAM_DQ;
output                      DRAM_LDQM;
output                      DRAM_UDQM;
output                      DRAM_RAS_N;
output                      DRAM_WE_N;




//=======================================================
//  REG/WIRE declarations
//=======================================================
// Input and output declarations
logic CLK_50M;
logic  [9:0] LED;
assign CLK_50M =  CLOCK_50;
assign LEDR[9:0] = LED[9:0];
wire reset;
assign reset =~KEY[3];

//Character definitions




//wire decleration
    
	 
	 /////////////////clock divider for sampling clock code here//////////////////////////
	   logic sampling_clk;
Clock_divider U1(
.clock_in(CLK_50M),
.reset(1'b0),               // Clock divider for 22KHz 
.DIVISOR(32'd1042),   //32'd4545
.clock_out(sampling_clk)
);
logic sampling_clk_edge;
	  /////////////////clock divider for sampling clock code here//////////////////////////
	  
	  

	 
/////////////////clock 7200Hz and 50MHz syncronization and edge detection //////////////////////////
	   
/*
asyncsig U9(
    .clk(CLK_50M),
    .async_sig(CLK_7200),  //synchronizer for clock 50 and clock 7200 from my HW 1
    .out_sync_sig(clk_7200_sync)
);*/

edge_detect_gate U7(
.clk50(CLK_50M),      //direct CHU edge detector implementation
.reset(1'b0),
.clkother(sampling_clk),
.edge_clk(sampling_clk_edge)
);
/////////////////clock 7200Hz and 50MHz syncronization and edge detection //////////////////////////


/////////////////Flash Control modules //////////////////////////
	 wire            flash_mem_read;
wire            flash_mem_waitrequest;
wire    [22:0]  flash_mem_address;
wire    [31:0]  flash_mem_readdata;
wire            flash_mem_readdatavalid;
wire    [3:0]   flash_mem_byteenable;
assign writedata_left = audio_data;
	assign writedata_right = audio_data;
	assign read = 1'b0;
	
	logic signed[15:0] audio_data;
	 assign audio_data = data_out;

	/////////////////Flash Control modules //////////////////////////
logic pause,start;
	
	flashfsm U8 (.CLK50MHZ(CLK_50M), 
		.CLK_sampling(sampling_clk_edge),
		.flash_mem_readdatavalid(flash_mem_readdatavalid), 
		.flash_mem_waitrequest(flash_mem_waitrequest), 
		.flash_mem_readdata(flash_mem_readdata),           // Flash controller is fed syncrhonized edge detected sampling clock
		.reset(reset),
		.pause(pause),
		.start(start),
		.flash_mem_read(flash_mem_read), 
		.flash_mem_byteenable(flash_mem_byteenable), 
		.data_out(data_out), 
		.flash_mem_address(flash_mem_address),
    .dataenable(write)
		
		);
	
	flash flash_inst (
		.clk_clk                 (CLK_50M),
		.reset_reset_n           (1'b1),
		.flash_mem_write         (1'b0),
		.flash_mem_burstcount    (1'b1),
		.flash_mem_waitrequest   (flash_mem_waitrequest),
		.flash_mem_read          (flash_mem_read),
		.flash_mem_address       (flash_mem_address),
		.flash_mem_writedata     (),
		.flash_mem_readdata      (flash_mem_readdata),
		.flash_mem_readdatavalid (flash_mem_readdatavalid),
		.flash_mem_byteenable    (flash_mem_byteenable)
	);
	wire flash_mem_write;
	wire [31:0] flash_mem_writedata;
	wire [5:0] flash_mem_burstcount;
				
	assign flash_mem_write = 1'b0;
	assign flash_mem_writedata = 32'b0;  //as stated in lab manual, set writes to 0
	assign flash_mem_burstcount = 6'b000001;
	 
	 
	
	 
	 
	 
	 
	 
	 
	 
/////////////////final project code here//////////////////////////









//=====================================================================================
//
//  Seven-Segment and speed control
//
//=====================================================================================

SevenSegmentDisplayDecoder U12(HEX0, inHEX0);
SevenSegmentDisplayDecoder U13(HEX1, inHEX1);
SevenSegmentDisplayDecoder U14(HEX2, inHEX2);
SevenSegmentDisplayDecoder U15(HEX3, inHEX3);
SevenSegmentDisplayDecoder U16(HEX4, inHEX4);
SevenSegmentDisplayDecoder U17(HEX5, inHEX5);
  logic [3:0]inHEX0;
  logic [3:0]inHEX1;
  logic [3:0]inHEX2;
  logic [3:0]inHEX3;
  logic [3:0]inHEX4;
  logic [3:0]inHEX5;
  /*assign inHEX0 = phoneme_sel[3:0];
  assign inHEX1 = phoneme_sel[7:4];
  assign inHEX2 =flash_mem_address[3:0];
  assign inHEX3 =flash_mem_address[7:4];
  assign inHEX4 = data_out[3:0];
  assign inHEX5 = data_out[7:4];
  */





/////////////////////////////////////////////////////////////////////////////////
// Audio CODEC interface. 
//
// The interface consists of the following wires:
// read_ready, write_ready - CODEC ready for read/write operation 
// readdata_left, readdata_right - left and right channel data from the CODEC
// read - send data from the CODEC (both channels)
// writedata_left, writedata_right - left and right channel data to the CODEC
// write - send data to the CODEC (both channels)
// AUD_* - should connect to top-level entity I/O of the same name.
//         These signals go directly to the Audio CODEC
// I2C_* - should connect to top-level entity I/O of the same name.
//         These signals go directly to the Audio/Video Config module
/////////////////////////////////////////////////////////////////////////////////
	clock_generator my_clock_gen(
		// inputs
		CLOCK2_50,
		reset,

		// outputs
		AUD_XCK
	);

	audio_and_video_config cfg(
		// Inputs
		CLOCK_50,
		reset,

		// Bidirectionals
		FPGA_I2C_SDAT,
		FPGA_I2C_SCLK
	);

	audio_codec codec(
		// Inputs
		CLOCK_50,
		reset,

		read,	write,
		writedata_left, writedata_right,

		AUD_ADCDAT,

		// Bidirectionals
		AUD_BCLK,
		AUD_ADCLRCK,
		AUD_DACLRCK,

		// Outputs
		read_ready, write_ready,
		readdata_left, readdata_right,
		AUD_DACDAT
	);

endmodule
