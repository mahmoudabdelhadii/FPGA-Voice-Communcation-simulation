��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��,�y�}�ǰ�=4d�H���`I"��W�`r���T:tB�T4D�m�)�	1��I�t��
��8(�8t>s)ו�."[�漆���]�~�]��;�O(1#5�-� 偙O��QZ��~rL'�x[�i,mׇp���O�I43��4d�,�H�����SN��d���3���r��m���̨T�I;uj2Y� Er�*p�Q$Gm���p�V�`�2^���,hz�<p��l�Bxt�5��s��\yq���#�@W���f:m��T�	,*�񞭋����_��㧋l�	�\�:��uGd��PǷ��N�I��_����Tuv� ���us�(H�~�{2H�:Zor�Q	#%�3ˠ!��iS��95�,?�.���/�F�i{#���Tp5����Ҥ0{%���2vpn���X�����@l����3dc�ק�3	�Ed&3�ZN O���z��s�yxӡt��v*}ԫy nj#��lc��m戭k[��5)�A#�����8�!�]�Z�s�M���t��w�!��'ÒE�rv��Ϝ�c@<U��\tq+��&|�&X1)C�����r�A~��B�&�����s�:n{p��͠R�X⺂L^��R����c���f��J^?��ܣR�O 1�rV���:��T�4���AD����˩�F�w��)Dm�O�b,�a���1$��c��7t[i2>�ޔ0,S���󧇳Ϟ�ᒨ�-��}�!6��Jyv�醊�^_�(�H�(y^����o#����X��3-�k\8�M�T�"`R�DF6ȕ� �,5�;Ҭ C�k���1\������k�t־9�}���� ���QHF��"��t�9 ?��{E_�7��!����](�S��0�q��w�9��=�i]�1�GʦȪc�W�XC�|�$��}q�6����zf(����լml�dz������*�eLD�*�,�m�]ہ6����D�Gw� �g��' A���FX��\өܹ&�6�h�Ð�$�(+��埧��= Eza ��찠pr[�c&��nP��x�2�TK�M�V���3Y4vIR\������ɭ�1՟?4�_y�y+����ƄJMm����@����m�����c�t�����:ud�Q�����T4���QxBŎ��\o���t�*Z�$�*7<�t~eP/`lfhg��6��[nn��#<����n�D:� ����4��y��I�I$�c�	ꈞ����G�l�\a��~�a-�]EA��|I�{��#�N�e�R�+Ø��fyz���%]��?��*��XGa{��!�N�\�$� �˨T9,B�-��Bt�S�Ft4�V�8n\)�Gc�B�b��5��]Y7�1��ȴ�OvG��Κ��ئ>�'�_��M����0��*?���$���aο�Ԙ��	e7!�
������3�>L�zcA���ฉQ�!8@�3nd�~����PU �`���1:�hr����+��S�w���"&�(��B/$��]T�ҢY)x�+��+��9eC!?�%)31�Q4����
@��� ��pz{%Q�$��ǿF���0~S�`L���;�����8W��u��:���#!4b�hn��JBl�	� ����:ӊ#�v��p7}`<��-���U�;���3���g���sG��-7Ԧ~�8���$;�X��&�}8|H=H
�O��X��W���b�mh�!���p�7����J�
�h��^Ly���Q+����?Z�2�jh��B��$��\�9+��|f+�f4��+�m;��×�o�����Xx �	�ۆ�,�ct���K~�"���Ob�P�~�B}8�*���{�Glj>
�c��[&�&���XV�#���}7;1�%�}�F�>O.	(��4y��d*9<���m�W�v�ō�ʱ�wj�W����=H1C{���4E�Q#�UB%ѣo��Q�rD���z�0@Ԇ�׎L	��	~�*���i��K6P��#I%��kD�d]��b�[��	j��k9����j�(uB���YX}v9}�18�l�k�Xg���(U����ϡ<->�%oe֖�L�!���H��`6]�Oc�yo$ ��`��y���癷��y�[ɟ��O�s6��h@�T�5]4�-�GS��$�b�Ě�����zY`��.MI��墟�H�d���� �(M�_�`�c�����>:n����@��V���-����a���Թ*��eQ6K�Ÿ��o�=��x}l'j��#�T$���lm߭V���8��z?`�I������q^	C]Z~YRvB�]b����L<v�U�n�y6\^*] _�-�I��.�qm)9Jt��Rk&��t�|���IY�U�˶I�y)XA�n7��I�5��D�u��$IL��|�$��,|��=s�.mD� ����*`|��P����	�7r?ŞM3�l�7��MA��lf�ܲ�yg���*��a�K_+%�2sE���=9> �<�J�� �YY� Z���W����D�DwL�wX�2����T4�w>��}�v��-��`lH���G6M��r���������/z�`0�#�G������9J�I�E&���:\@dm��Yi���"�<W>([C�-��Kȶ�C���!#�b�k̏H����p�d	2���hE�7�w��?���#��n�D�Wڵ^4L���P(w�٣���J���|���?����X [�E�����`R�f�q������l߱p<7��u5��<x2���� ~*��:�||��U͒���?ؓtT-�:p|@���Y؄���ؗM���"s��Hŷ����e���9/N��n���eܢ�V_y�����TA=�jж�SF�1�Nl;�uOҾ�l��*�O�V.���W0�F9�����.`ۣ��Vܼ��0Ob#y���1ad�qf���l��=~�\=9H��3ф5�Ҿ���Z-��������JT���#������#s調�<�����:V�I�t :���IV����9�р�Pm�`?o��9;��S��5��K�}��\�G�����)�:�M5��"�C�Q;Rn��
(��2�B��,��"��D'��P�B�X��O�"��a̞�4�e�X8�Fm��B����@����ތ��EC�vE��B3�����A?�H�;V�~�R����Ę���'�٬prYz��E4#�V���L�j�XV��X^��
�r;�U�2-��1�tv�������H�i%��m�=G��D�#t_Ṕ�~��E@�a���U{$n!�(��*�)����S�?f�_u�#����M����>�>J� j��#O�w��y�$< ����5 3kS��f���}���iU����B��i�ҍ