// RSdecoder.v

// Generated using ACDS version 16.1 196

`timescale 1 ps / 1 ps
module RSdecoder (
		input  wire        clk_clk,         //   clk.clk
		input  wire        in_valid,        //    in.valid
		input  wire [79:0] in_symbols_in,   //      .symbols_in
		output wire        out_valid,       //   out.valid
		output wire [4:0]  out_errors_out,  //      .errors_out
		output wire [0:0]  out_decfail,     //      .decfail
		output wire [79:0] out_symbols_out, //      .symbols_out
		input  wire        reset_reset_n    // reset.reset_n
	);

	RSdecoder_highspeed_rs_0 #(
		.CHANNEL        (1),
		.BITSPERSYMBOL  (8),
		.N              (255),
		.IRRPOL         (285),
		.PAR            (10),
		.BMSPEED        (1),
		.USERAM         (1),
		.USETRUEDUALRAM (1),
		.USEECCFORRAM   (0),
		.USE_BKP        (0),
		.USE_BYPASS     (0)
	) highspeed_rs_0 (
		.clk_clk         (clk_clk),         //   clk.clk
		.reset_reset_n   (reset_reset_n),   // reset.reset_n
		.in_valid        (in_valid),        //    in.valid
		.in_symbols_in   (in_symbols_in),   //      .symbols_in
		.out_valid       (out_valid),       //   out.valid
		.out_errors_out  (out_errors_out),  //      .errors_out
		.out_decfail     (out_decfail),     //      .decfail
		.out_symbols_out (out_symbols_out)  //      .symbols_out
	);

endmodule
