��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����N~@#�k�0!����+��=L���0�ԴZ�2�Mc���ZO�����=�����վ�	"cqw��a��TS[��{=:�����K��-�մ�(��k��N�-� 偙O��QZ��~rL'�x[�i,mׇp���O�I43��4d�,�H�����SN��d���3���r��m���̨T�I;uj2Y� Er�*p�Q$Gm���p�V�`�2^���,hz�<p��l�Bxt�5��s��\yq���#�@W���f:m��T�	,*�񞭋����_��㧋l�	�\�:��uGd��PǷ��N�I��_����Tuv� ���us�(H�~�{2H�:Zor�Q	#%�3ˠ!��iS��95�,?�.���/�F�i{#���Tp5����Ҥ0{%���2vpn���X�����@l����3dc�ק�3	�Ed&3�ZN O���z��s�yxӡt��v*}ԫy nj#��lc��m戭k[��5)�A#�����8�!�]�Z�s�M���t��w�!��'ÒE�rv��Ϝ�c@<U��\tq+��&|�&X1)C�����r�A~��B�&�����s�:n{p��͠R�X⺂L^��R����c���f��J^?��ܣR�O 1�rV���:��T�4���AD����˩�F�w��)Dm�O�b,�a���1$��c��7t[i2>�ޔ0,S���󧇳Ϟ�ᒨ�-��}�!6��Jyv�醊�^_�(�H�(y^����o#����X��3-�k\8�M�T�"`R�DF6ȕ� �,5�;Ҭ C�k���1\������k�t־9�}���� ���QHF��"��t�9 ?��{E_�7��!����]k�j*�Q��~�=�0z����o<���_TC?�];iW��M������O���R�$�lIlqֿT����N�B���ڊΑ��R���s5��yEK@aTaz�]���@	Ɔ������)ɏ�������7~v��ROf��!wg��K,���Ҭ�#oВ��/�~�+�Xp��k5�����	g4Fड़�Sw��%���f���H����]�e-�I��-$�;5����r��� ,*�	D����CE߈H���cBIh�5!���v�Gj	�f%<�g��d� s����YßM�����KA�uV�,�B��(��BkF���ڮ������M\J���cr���C?��r��!���F]ad���&�~�%���;�VDko	oB��>	�����.��S�L�$�ݣ���fj��e&Qjq������a�A�V��]R��·\�J�@��z�8!���n�͊܇����K��#yh��,jƆT5�m��^��*F:�*u2�������3�C7� /�4Nb(A<�� _�@�b�}��v���R��E8�,��:¨C?�yl�҅݌u�A(�+~F{Y�D��ch���d��&x�-$Y��:��ז�ś����N�#�J�~1�w�.�k� ��V�{�h �KzФXy뺿E��-P��icUNZ��) �hR�������������LB3
k�X�������ʁ'�����ѯ��1�^�LerBZ�#-������߮� 
�Ǔ����A{NBIbS��K�0H����M��3�Nu��KY�g~̦
�������)��2�����(ĻD�"�ฎ7�->����B�2���Sq��^l���_׫�p�����r+�a�=D�s���(K\�X��^&��Τ�[��F;&܃��BrZ��؛��Y�,\c	S}��������9�@
��M
����˳�ee���:��,��SȬ��4��� �;g
�<�٣N�];���%�y��O���.���S�!��x��?�H��G�����_>�Tc������a��f�/6^k�v�-t��+��#l��p˙���G ��K��	��9*�!1�����>�{�ഗ�iQ���ܯ�)��������"� &�G쩰1].2��Z,��-V��h��)	��n�\��Qm���g6�^=! �yS>a� 5�Ɋh�����ݚ&{�9_�{�Pl�eܳ�R�z�d���f�Sװō���bs�T��(jxBݸ?�	r��CͰbk���k{9�$���8"��Y���?!DC�|��ӱ���+�:�I�c������w�,*Z
��V��KaoN�7�&6K�(O"����Hܣ�fq���䀋���;�����`�O=^	��))`N"ao��՝�V�>�[-�l���L?�RPP�4{5ݝ��ݤNL��ˎL.�W���T�gl<�=HL��|w ��_F�3�4�WL^$�uHۼʏ��E,g��]��}O�wP���S�؊�۝L�&��/��/<cy$����	��0�b��Z:3ic��B���q��2��.r4��^�=�'^�#o3�Q��V
�,��q���b�p��Ԃ�:v���F�i���i4W�5G+}e"C��{��Քދ@Q�m\�`|M�A�%L��0|�۝�e�|�o�re�!r�}�	�� D�5.��!>1󆇝*R���i�n�3`{��<t��o�<L�s��b?0� �����T*�XҤ[�¬����Z���F�	��
�4�ݛO���փ,3��r0s/H�O��x�O�'��	u]K�܊�Mr�e���(��.�1�Y[ݺ�<\r0r!�����+���gu�%����X�E�pi����xN�4�$���j,�<*=M�_睹�^�2fSՠ��&.<��sWk]W����<�� ߽���I�a9n��1	=nppKR�mj����*�cO_1�@�JTr�p��@o���r�6$)��0-��#�qv���X=�y���C{_��e�Xx�@rm����I.���H�V�G�N�[
��e�.+��c����2�#��� 7V��OL��\/���cR���^k;f�̻R�wI�ŕ!Sa��H�WI�,�:�5�9('�FL�)�^�M�0��#�������<7�r����b�\T`|��9��u;��C�g��Br�!�J��~�.�7�ߊ�&�{PڟG�w'̀���M�u4s���o��\=ժ��2�h�k0��x5w�}?�lBQ��Qф��"��L�����I��T�j�l�0}�ya[����~�F���\�3�ƣtg��N�
m=�:��ӽ"d?Q���"+���G�R}���s�CbgM��
����9���^>��=�ύ�8Ew��";D�L�>��(��]���:='�B�hwEń/���29�X�{u��P�ij>�jQ�� ��[^1�w��<�@�Թ���&|[9�_1�Ϋ�_�d;���E�cz�/oP���֢��v�����Ұ��/�+�����t��:q���垡zV���4nY�R��\�:��3kϹ���C:�(�s��""}cG�>�8�?r��y1 N��^
�[7tj�����y=Ԡ�`�P��2�KB)��׷w��|�e�$��q%��+�����M��ժ�c�Y��tp)s9:��>O0g'���rs�O;�n�^'�����m�t ��8�ְ ���r;F]*ʑn�
��E訍j$�n��ΩtKB��C�~��s���mX��~��=Ts����%���߭cm1�0��&g'�`��-
�
��.!$��qրʯ\���:1w�~#=Ӟ=�+��ln�$�I�T��v<oA"��#"+��*��ܛ�U�.����LZ}B�����J`�1B�UT]\��d�,��v5!ɳM�Ss� E�zL�l��O��tjmZu$1Y�J��0�7^�U����LJI5c���\�hz����J����ה��K~G�g?�܎�J1U��?��N�Z 0+򙯎�S�JDM�j�7ؗbх8-J�� mSu3d��L����|��3�]�{�%�AEn��3Y�P�\2����[�]�,}�OcU���>��	N�c�%r��:�s��Ua�������!T�(^��.1p�f�X�u3+[cks�������O���7�I%�n�,�La'���!Z�´W�U{�,�تUV3!�'6An}Ǌ�7���LT�]T�/aö�(l^|��'L��R��Y�Y�.���(��GWE��Fn�V�D�J�ۺ_O܊��QLd��H-ٿ���{C�>�~B�֓O�+b��>�F��Ǒ7�ht���=�Y�P��9�HEݶ��{r��b���u�.^]�r���VLNR�2[B���6F*��ݹ�����f0c���j���F�������(���'�h��l��3v�F��Q�2]ǲ�<|=^&�F�\��O		��|'l:��B]��	�]w���T�h��"ݖ��F���u~x^���������>xM�%��ڀ�X�K��}k���1�?�%b⊣x"��CA����n�4�\m!�J6��^8�$�K`��3���.�[������dx�=e�v��G��ʍb���]�(��O�'F��O���L-3�GN�� p���F)��e�2�  R�z����<�i��oe�V��`Z��ծT����~]*����:=vR�Åy�S&Z�J�����_|�HP�ū{m�Q����×:tw��P�(_P��[�I�N�g:m���A*߉�A���"y'(��=��x�3�C]$�w��lT�'�	���ܳ�T`��+���]Ӯ���IW���A�c�H>��<I!���Ӕ=mP��uR���Q�؋zp����+ކ��,�۔�I�[��/�Z�����9�M����1��;��k=5S7#D���0�hafQ�T&6#���	ds ඏ
�����Y�:4���U4�p���=��P����)�q�J o�qJ�X쳆̆�&捓��k~v��d����M{����5֏F���⦵��� ��% k��L�!��q��)��!��p��d�8�O�P�O��.!p����o�'����Nm�ç��|u�kwak�lU�ۖ	MУW�>�HJj&HZ�"`��XB0AGU�֡����ɸ�ӎV[�Þ�Py�B�{{�T���5C�b�0p������ʚHL̑�Bx�b�����6[x�?�f���&�]x�c�w��ߣ���1�|� XK�nջ؈Q�t�B%k>V=��w�G�յO'�����u:Z_p�-�aC��������%29YJpo���1\^a�8%��� Q��$�~~;Sw��֟S�#�\��QwX�<y��2BU�W�p�# �Gj
S�M��U�1���f�G�;|P�!�?����ҍl��A��T4r`x�s��o���w�Ր�3���h�É�4�&g��_�3�N��IC�l�Z7�:����N�E-�xu��T���a�`����9s���܁H���kg�]L�]�]��ʖC]j�CI�Í������e�P#����P2*R����i]�IIu�eT;GS �4�����7l~yj�S~C��@������4���K�8���86�Ïi��H���lL�4~FC�����y!r�XucF�*b\�!�+۰5��ƨ��6eӜ2i���80�Vd���X�od2ZU��A(��?=��7��bXܢ�R����t#�(�l_o1T(^���~1���Q�.�Ɵ���6�\�Q,5E2�%��?��y
�Ia!�R\*KL�8J��|Ȕ�(z�`�����f�\cm9��RR�e�6`>z�e�)��h)_��x����><�F5�p��z��W\&8��^?�����x�g���֙��E� uv�6G)�w �!`
\�gC��+K]cFt�WDd[T�R���d$�'�����;�#��?⍘�G*>м�&����~aE��$�ˢ���xQ�YI�|<?:��R2�_���߭X�,�3'}�mn�4*=c�{?�*�?r\�+���W��V9�˖Ft��ms3b�c�U7�C��d4@�F�L)��H8�;�wf�}��L�7�d	��~��%���sg�<���!��t����z_o�u�)�K�3���c%W���1�A7��d��|����|�(4:s����'�{����� %w� �֝�.�-�3�^!-궄R}��))�3�W��;�|��9��yG���L��%��r��RC�3x'1���Z�����)%o����I�e"iq�'��/a�����a���Hq�
�����1�̿*��ٰd��bk���4�c�%��x����!
R����՚nˠuq5z��J+>�.ƪqk���g<��p���Y�#ȑ}H�YA�BET��H ����/�� �2��,�}X�d�y�@�`\������C֑��
�5��b V]er��3��H�|�vZO�inv��f��g��1�B��9�]�*�f���?���p�m�ڡZ�U�;��=��ׇ��8�)f�$�����aJ�~��p"��^b��F/a&ڦft�ܟ��/�T��4*�����-ĕ�8��l��t�Gf]%F�,|iB���E��1'A���I��r+� z-���0ԩ:	I�PUE���ӟ`��QpB$VN��>���(e2�	�`@<ʗ�-��g_�S�!�0X�s6
}T�}|ZfP�]��G1�1ֵ�=i�6@��)	'$@~'�=�5aJ��]�)�O����|z�k�~��2����5����MX#v�.L�ɴ��Bς@�I��6J�᜼��n �1^h:Bt�:z&�i��� 0�B~�¹�j�p�F���H���[�
q(+z�й�k�˸f1�8�&w.Jh�Q��)¬_�ӹ];�R�P�����]j��*����5�{rՃǬ����(@Qd��6�qG��&jn3h���m�+����nn��)L�Y$0��>��t�d��5k���Zz_�D�T�'t}tZ��I�T�d0Hf�p�a��.2���>��O��J�W���
���D��-�]s5;$�^�K��� ��2��65�Űl���#�����܂�!�C*��e�6�}���?�S+n��-Pu�1�s������gI�c�ѳ�{�;꥔p	X���>Iu�
>���#>ǘ�/u�I4=�kS	L���Y�8M���A!����ְ%�AZy��
�$Dʾ�`�����ԗ���<���LQb.}�Բ���#�꾶Gh4-��}qξ��ڎO�Ǯ�Lk� �	�$
�k �5<"�N���h%��<��ʬ�0I�T�R܃��D,�A��x(���"@�@T��a�O�`"�i��Ĵ��'ypth�(!/����=8�+��Dr����4�n��E+�|c��AL�ŖD��$�Y�7�?��/f�Q��������<�Z�]��ʾ|���2X��e�%�8�Ո5�?~�G��5��$	��A�Ʉ-���-h���)�7az:z�wŢ&!��� �&>��'�f�@Il$�������#U/1����zFj�`P�,��S�O���7�S�W୕?��M�H�Ԗn�&C<q9���C�<!�����jZ?�ո����N���;�R�亂T�1�������$6f�e�%��2�ĝc�����w�L~��9��\��1�y*���L`��H+�i��Q�W�>�4@�N�Z@�F�v-��^�j��wlx�Tq�;��Ssf���'�	�m�����~��6�G^����	�+��2E���奡�\����O��D"(H*Cu�)�����M����NlD����K��4�收�nV���VFFq�=$�&�f���?H#�{�*��}�埑������M� +��̿����5�F�M��x�'�?�aa���όgx��!r��>�^2����3�������{2�;��T_r�(m��6�]"O���|9���v[�$�L�I�T�fӞ.�%,W���xP�1W�+��.cd����r^�6yp�XVV�{&T��C��*I��BP�d�]^]qk�9R���R��^�G��ξ�B/�o�\��1��a���Kg�R�ȕ�l'��k�	�u��:i��Yo�?����ع[�_;� �gA�@��J��|����U~�K)��p���V�t�n�gR;n�#�`
�-�
��OZ7��wzN�
�x��2N���1!b꨸�Uw,��gR�ESa���A���6B)�]�U�}��1������w�slqߑ2�1|A��጗ԙ2�;	��Х����!�8Y����ɽu�"��
�2��eN�,����p��s�M�����|�Ug�v�9��yJ���t�MR���  
�a��O� ���4�%{�+x����9IW�
8y��j�*������^���������-�Xpı}�"m�� �:�=�/wb��8��1Z��o6l�'�D+0��E�J��蓢�41�����]Ey%5�]�wD��]����`��G軧��\���k ֑j9���[����ˏX���ì�d�n���l���Q[��4oj����חX�K9Ot� )X�7-�m����$8�IxW� �`)�g���"Yb���>�"�L��E�@
"7�x��a�zdi{�B��.BJ��t���y~��������KZr��6$��[kri�|�JR���KV�*fw�(@��͙H��Z션&��{���~�i�b�	 �@^�� �&�'�00����HTB��>D�m	Y�[�����_���Xq^&_�q%�Vz7�$0�������"�i��!�搯��&(D�f\�W��YeVKvV�6����`V�dk�3=/N��Np3�0|�w�ҧ����r�f-�?�Ԥ�B/�P�	�O �(���{/ɶ;�k����Wty�F�uMb����O�<=8��~�� ��8���k�%�-�I�����9�aΔ�E'!�W����~"�|U���K��h^ְ�X�p�wd Ф\5�`	
�N�ke�٬�H62��gb:�.��W��oAnn ��̿�����sJH�W���<d�Wi�ɖ��Jq㴪�#F��a)���Q�tR	|���Ĭj�@S}��>qZU b�No��a;0�������2���!I��%6����mj4FM��zu"��oԽ��nR��ac��3c�04
����2Y�0�:U]�^�*����H	�a�j��bt�9�:"�;��$M��
E�VÄ6��n��Wx:�5)����kk�gx_��X,N7��5/����U،�~5���}�ikٽ(ēo<�?=�	��kyh����XtT���ŲS����=�Ҽ&�S�
kZ'���n?���r\����]�VEP����}��S�@C�;�V,�)A��۫����O5�Zoi�5�NC����԰����_��Ah�5�E�oP`v?�ӗ,���N¸=��;&r�y�sxv>A�>�s��՛��I��� �O`����C4����߇1�i��7��
VӖ;�k ��Ub����t�=�����իp��7����4�O�0��;ƁO�C��R� ��ſ*���L�R�Wd��KV�遴��B��������ެ�罘#M��Q�}�(��C���T����q{U]V���E�Pⱶ�6�k�u�~ϭW�4�&��@9Zv�������hD�[(a�j�m�Ͽ	�.�S㐎�l��ht���X(�3�Z�q ۣT�^���G"�TW�����Cr�II]a*���i/�4k�س�h~���:�B΢��x5��R/�Q�o0�ܨ�S�k{���[7f��ՒU�_�,�EP���9U!Z[J�"G�Ԝ�B`�k�/�w�P�'捥}q�a������`�S@9{�gK� ��W�ݴ`6���d�p�d�Gft���ȱ1A�杄�K���� ��No9D�NǉO�>���{:�׏)��pl�R�Q��[?bN�;�y�����)�
Tϝ���rMm�p\�e=pLG����8^���obg��/�К}܋����Tv��!R��
�bS���3^aM����ݥ��}���q�?+�X0�G�ʶ��櫯�.@�?"���A��Z'V�M���Ċ#����+o�riP:T�0��Q���ZX	�ndl	�}�o��[�����T��@���`pb��w�xo�He��D$��� ˓�����K}���-H�dB�+?�y9��{�jP�t�7��y� [���R4�����pB~����:�0�c���� ��@��\�j��r(z��T!�e���k����	~v�s��"G��֐� ܶ�UY7��X����C���ơ���o�h|2����0�pN^�X����;:���N?�+�=�k�������F�󉭯�IX��r���}��m��[$i����2WΓG��d���d�%T�$5^z+�&�W` 1IQN�T�ᛊLpg=�&���~w���bA�J�(�A�X!w�p��d�m6������?�AQ��F� (�a��foI2F#�Gh�-$�����Ɯ��\CG��;/�r͖.4�))æ2�J�e��~�ظk����_�����,�̹�py�p�z�šH��QW3�]�s�{���ɡ(O��s��&����õK�[^�9_�����E��^44C��1U�Iqz)��μ�uR�ĉO�J)��|4DS,=��"-��q�{��\�c(�OYYM�>�"���Lq�hm���]�<IGӧ�7�n��r�g�x�I��6�ʎg��z��A//�}|	���L�\�ַ��1�
�,Ѷt���Z����wM3p�:P[�ڶ3� 1�΢�'*����_Tk0{~k��W}�2���l���؊q�F�9�f�v)z^���>��!8[�nF�4���;�V?]�Ca��1��f���ԧ��wv��m$!n
�S7�
����i�+�'Xհ�{�G��(}Bb�(�v��F�Bl���}��f	T��mt��|�6d?!m y���o�/øϸwJ���J1��07�z2�酧2 ��`��"kTN��+'(�L�d2�%��S&��G$(�����T����~�j'��ψ�X@��a�A��P���0����I>��S~�$Lh1�lFY�/s+q���#$o�Gm�G(A3���`�7OX�3|Lq1�7>[����� r�����&��
�����JBV2�0�^���(r~&��5?M�l3��T�m��7� 0�@�w��~���'xsV���͎׼KSh��%8/.���T�ek%�x�g��yOl���+|�������q��e���eIT��?
1L����A�b��Z4�C1kƒ*�� �5��� rȭf�z�ٸ1����� ��|o�\�
'R�#�-����M��-^��j�h'����o��j'���l1��
���梏2�q���*��C�
�1$b����o��1
�Qqf�-Ok)c�hMBy��#����i*�>�pt����������Q�3�5]uYX��ʫl��(�s�k�V��cϻ��_g6�rn_�����Q�Z����^=.��ڜ_J���.ȉ)���� 1쮠(����{�I�9]S`�.}Sx�6�ȗ5!p��J�D ��0�z�%�oRT��y3���;yu;�+���d�(/�������揦��X��p>�� +b�"�e�&���M��7��6�@d��S�_�+��p�R��V�G<�"�Y����?9t�q��t�d�m�Α��p�5:ȗ��������B궃 uT����І{�6G_l	�@�7�7�j9��[�e�K�q��:�1�R;��'TЁ��WH�N\"��"��t��}7��s���<ӳI�Yی��4��[ۺ�| �H�G[%��hDѵ���X���tr�n��Q|���w��Z�Q�\�����Cxl�m�e�����|��v��,ٓ�\{JQ5��Nv0��Մm�̋,�ȠP�ĭ!���.]�!�զEq���}��Sx��:��o��@c���*�i��Ԇp��=�8��C]jq��2���7vG�������O�o凮��������q�v����R�ը_
֟�0m.��dn��A;�B� �u0O��1)����G��~��
�Ε�K�u���o�朽 n.y�x`��|���8����SñK�]9���