-- (C) 2001-2016 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
vcU/Sp1RgXbOpR7yavQDZCtrAypB4z1bU323X32jkZtR5RYUmS88rRe68QKatfRwbQ7ky5WQn0oS
KyY3kDGNssYgWJUX4B/L1cZR68GSNEeJkFdFTq6p9ofVFOo/zA3ZtHqPuFrh+whuOtwfcW74TCXt
AATVv4jidg0XhvJzfUdfXReRSMkhQdhWDFPyIUhfd6xCPmUlQiB0I+SgusQs9KjAnxHoO8JjdP1q
/2z4zU8ieTMTyInLgwKOnneC6NepptLhu57Bkyg+GIuoJjB1MtzgWmjHSGkwdRnxl9m3hfoeB5Ux
lavqDx4IX6Efb7pTwKZQ5DEks19vGw90FRW6pg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 2336)
`protect data_block
JgbEhYciHgt3olunEyxejA8DULt84ZrqL0qrg5vSH9TdMp/z2/b86c5W4V9yGnhgBR3KAIG7az35
6imx9R2ChSnPyKG2s3tyYbM1BjVhjW5e8221tgIDgvJTWR9zf8LiZDMKwKJW//blc+VVT+SQWfx2
VlYk8bOa3E9RTt8Fv9Gv/46Ca210MTSYeGw0wQqYAJJMj/OS9wPToWa/igh5mC8k+MGfSQJw+ojF
vOKpBpml29N/Q8XKAA/yXz9Fx443uyFtTAcyzf2HK+bFO8bl4Ds8C8zAQWdwXFbqxsc3afHCYEut
3J2s68WQAW59G0w1L0HWLqBqA2UaTYLWYLbYI1qJ0etmf/Z5Jvukdt/tKov+TA5vxJIEL7y2NCWB
Foj2r0KWZFsejwNuRz5nHslaGVltV9grQbErP+NGex4O44pUQUqknRiKHMYHxtNBHR5cjPe2GeVZ
rzLVTm8pl9xIMONb1ep/F5+6S8yTO9wVwk1oBOGAITg+NlfAUAc+1TSLOHdF1XKSFQIUs/KdGb9h
c73u75RtF0dUpKpn2sIMAxGJhG5t1ZQ6senzg/9uL2/P68HQSRbXzl4gS9J27ITGvMSPXMwoMV9i
c10xZR0OrfDhjTOR4O/6uKJqJrJSSal65yFojaN8qOCPBhHuNGKR+HcivXcIWBtW+rxXNmC8qlTp
lsE0GX/ZVCvaN1MYTPHeZvLJtPtXL2epa2QQGNwFQGTVCTQspjFVQPewpTAPn/8S3RW5V7FqTPt8
yu9uHFmHRaZ4ErvvZpVpE1DJkvpnF84YMcbtsu2s40g5qmLYXmrEluQ5GilxOAnBKjs8VY1DCoXa
6Il2FeF7gtY23RZP4nWywbyq0rVmvAjm6Sic14JMtnKbGi2iDSAciMlGaAY28CS/XdYYUpjf3BpL
Ec6LxK7C91gNDYXbIQhGbCIbYp3atw2uzz1YYdV+o99KeQuQYcZXvMQbSIoOhgWMcHs5DsqovZI5
Kny29YED1tiI8l76NQhVTDPs+c1pa6mLDV0fwv14yTcPvRaQNZVwGH5zGIVpC+0zTfnCQoDdli8X
UWnHML2z239g4mpjnigOgq/CD0EUVUjOM8Hw++fnk8DUyvCyPzI6hUlzRsnueP5Uaj5e0uA+kymp
zhWK9wHe/QCkSkik2DXHzkG5YieIK/6NF2GTq4YfyYwHiCYZJpIPsqD3AhO/NhP00cAAM9EguS+4
yAWmebnFrl6ttov5sC6MTFVwZITuG4wURmpAVbZk3ElpXmCGV9sqSe+fs4gH58PHcSi8SDuScbcZ
4yblofJFvocjiFmL7TFcoEYUJSy1rUKkIcnb7DX9JgIwI65zWMGz/djLp9VTs9w2zr8ey+2TcRpB
487zHhp+GeNOIuY0aMZYwO5x1ui1Sd//3HB4xfd3+Oh6mvbU7evgSQx3hhPU3b6Q9BwarfrIgDrC
vW00K4bpOQXiTmnPcawxWRc5nnwzQHs0Bfx/UmGMeQAlNPkTd8nGtaUg9M1cZixHp1lyXhu35CTO
lVf+8PlEDKUAAkQ7EJXYT6IR0MHM+Ae2qySs7f5Ie/gktWaxhuAWQJtprR/l9aocRVRQwbE9JZJ+
vk8tRmfKMR3vtmeQ4pG9wbi3YsJR91q2q3Nzu6Ljcj3U8gMOUJC05sfWt5dI+Xs0ZflLtYbyfAQV
oUz6alSNYi952E70qTsuqONq5ilwys87VBgNkElNosMJI656kLmZ1D0iMVhhjcdPQOnZy6fAw6W9
EJxwSAiKbAzwA9ece8JT607w81TQrwc7I2wa7AqRrhqnWXFgRu0KCctDnptbASyE2ILMCIG2fVyt
+j9rtX3+SAQwHHOBSRE/f2ZKRbdOveXFsqPL6A5viMx8ARLCR3Ta41/RN1h5C7eNOuBNRuC4Udg5
L3qgBYcuJrbibIeL8I2/02lxBI5RUyinpH1ip4t2aNvbbdzTt56zpXbT1qp1vgiDebfkzykBNEk0
FPTDYCDpVTIUGYEKxd8uZohNDXBiloruJzeJw0kzEnFWEgZ8C2PXZN4ZFGliCPysuIPRpfl6Wv5O
0rPw80Kosz7ydmq7HBVN7b5fHlSBThMYryN9aQbzd8u6pccvTqBtjFMl2z99Lun5L9donu9H1URX
rrQ4FtAFOKy+0B7+NWZm8+PJsuEYN2jAwoASX4mMUnJB7lotY8SXs7OTS6cjlBYHdabUbTCavNZi
VyrKZww6ip889wWsXTpc3sDbAUWKy3AobNkfyD0pfWhqEEnem/2gzXhnwqSbPDujyk5X2Ui4YYRw
/vch8d3XBlSpxhYhbXAUujXBeQHdWyeGBsjNoq5OospF3VcF9dDYE5l4r4B52ICeNARMtpeIQ/h6
4YJHnTl1uhaBoAmmwTGH2VMKv8vu4cN2ekYhQuqsos+mCexBzZd4r06V6P2PDqKsw7trJwUpJxzU
SXaSIlgdWsZG39RPdMxxAdnlp0xaSLWE8EqdnFKPwU72st3phdOAE/Ir7G+hhnvvoB8YrePXUi2w
5+5bVe2MeROMVufeM6Ww0FiTcpFlt4wdZQpGo8iHxGEFu2h+Uawqs7nVXWvDsKh4QQktfg5FhgW3
bHFQu4avYIEvKtjbShkmLS99Ek3xql8CrtAX0BoTzeZduFD5k1+qPsEIMWxH4MhocEblJ4dvoao5
zhAK7lWThHKP0jxceDYLnigxKxYU7uiiTuHPhKz7BTGdhFZBGjKPyF/HXsPq1WyjomEbfOdb4nxe
sA6G9phAizuTYd+MyoAdh4qlAI9/gWsCgaKzUF5kf2vZc8HdX+WP8N2ZpOeG9f1cajjrhPlCdgtS
/bZNi9TJrRo6p7MrDdC7Rp9H7yHFMkiSxZHct1yZ+PlRpiKF3OjJlGeuY5QF80/jwyCac/Xh7g9Q
mS1lyV2xmZwG1v18xR3ti6c0Yie7jfbLqTHs4WbY/c/IKfKVD+tjvDs55PpKeQC4tfsE3yiL5zkH
bunkPu9e/f3XQHn0kRWW1HLmdqS6lHEicUtej7+z29pFJ8x8BWIPb05oLuq7C4Sdd+b7MXf7A4N/
oMYaG/yF+ZcfCX9cm4VAO9c3wnmeKOOXHSeDxyuXx4updU4GVI0jvrdq1GqThOPID+ovYgIvaJw=
`protect end_protected
