-- (C) 2001-2016 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
hq+hTK2Sw+8Iff4yoGmZv7N8g3EkUHXe47QSiz3vwbv5fMFVq1ATebdOr6J3H1cMO/yGBB1r8YOh
lvlnNoLwRFsiAdvdnX5RJL2bOw5wmNhUXm4vpFISzeajgf4pUAOhjuQqBBw6mZcBn2lsaC3UvrRe
FRhTpOal0LgSXmcIO8u6dsiAWyvbvq0Me0giDqeI91kHyXrGt4iK8t4eIAezFYXQn5sfIYVdlL7E
Goi9NkqKKj4zaGn2AkuMStZPjgE+LtkGz2/jrT0HsBy6o2oWR/+9E+djm6tkxWCrcj7On58vVMgv
lXno65nsNO5y0TTJsedOtjIRteR+zg5FVqHIUw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 26320)
`protect data_block
nNqSLa6XDrduBSCZC9lhwsSwvPsgeU8Rbo5m5oK3TJXAGm3LxF9272qbqMsevmEM/PqOsg4CSZij
TpNStcyzms83xlbnuENGb7GoLeTeuq9iyWnNE3SIzKXKoQfo7UHUOAK3dqUvWmumAtJwtXyMf23N
4e33+ZZNsV5UZrWEJyHuMtnxAKX/qCpNqzW8qTcnMfTG3NICHXj5GN19yVFvmpBm11wcvd+wy6IW
YD+NHy/DOAEVVC2CN/shyD6MGs44/TKzOwIMy8ROSofEc76/sRiLRO2OdANyRzTRc0ev/ows98wd
w0okKuRvq+eDl4bRO3AlFG4TYDU2KhG1llAydo19eiD9+asGhGGclI75trfaSOu2rXxNemZNtqo0
NZSrf5sUY7iyf/V6wqCQVA3ORujmrhOFP+9hge+BiK8XdslGFxke18jJ1Mlq4UqbhqBxLyfo2phM
C8WDmlmCwzrtId51z7Qau/0u74vVH6dGMpC25FdVN/GCzsO+mQuRe5aC0ny0jfDNX0F3L+J9bhOr
Q4hNNLJBaF8tnlG08hVY+6xIsLeBBZH5y0k+rXEQpcoCFO2TGWck9lTxwj+FAdEImjmpdctOxpng
rZ7j9805jkxBANIzXzeRwgLX8ZVM8+XmzJnmTaQ3UHIxE/BevSaSrGNunTGh9Az92XH6ZK6QM8M6
x/4pfUcBaPGoYuUQ5svEhdKb/OOxTl/AiLNjIOgFkm4AWlsXB1t/IkpQqvigbHYnCXZvOlEmAAfQ
hpsnzTMHQ0LYFjSDIfwXIGPuhBMdIE2NZB3WK1tiuBCfg41J0r2ZQGtyc7RMITpDmyQdR6dOb1LZ
6bka0ED93RsOZLVUklbLQaS+5TzFtYbCniit7frMrtx1JqiQZMSo9EzkM/wROrXQPForPDxGXpjw
1325L4LtPqHTRIyvBg1EVzSWg3iBU0neBjmaIFLUUtg4N6m2z4NBhjBysUlVAiC+FEDSC7xlDT9t
+dEH4Im2P+UrifZ3VZz7r6Av3wdmHxyRuvTcN87D744biQ/xQ/xABm4NTsQXX+fDd1El/QiuFYYi
1DSlgBCrmyN2NnmwHkkWpilVCAK6QQp1b3K5LZeZJKGBFSlgczZHAkRyyYBTioRaB/2X2b4Ws0II
PE0qs1dcVVZi3+dNw4LnR8NeXtV+OVaEMT29ohlPq74LStycKqMz1o81rIfeLR5c/zIHPjofOTd3
RkK1E5sSCbQgihwAnueE4t5Zvvp/t1gUWR+6WTeJGqnUVF+ynajDEAqbv931tzyQ7/cbvCfgjN9N
R+Se97k002ZuUzKDOeCV0P4aI3cKd6EYfSfJCZzJ3fp7KjfCpb+kynmcA7HVwwQHKg8PUFjSsST0
absth5NYMylJZWKf7stMswIK05gUathQPFclL/fzSJN64llUwmw6de0fpnlzbdq2Bx72/mXUDGEY
je23VdF51p5aVnbV4WAhDogz7lEaYuWCIt+QUM0fLClquiS5/4ZXZPuGSAdosH4ukH3v6QsFo9TP
WG97ECH6l6oMUvVvuXiBGG9goDnqqvE1Mly/4VSlDEvZz6cze/TYlnlnn/WiAoHeHjD1jRGWUKvi
1g2EdjHekom8CjkTnZgjBvX+n6GjWHVTBdppaG23Urxh2z7lZ93wd7Ig98qICNImETq0o+AamYAC
SKoUsiYi6TgoXmkn2h5GmUC9WGZQwoFAHbioayiOYUmpRhN3LYNDzKpY5fTTkE1EepqRm1PtHyvx
raKG70/ZlhVKE+EJOFD/Y3UevlTDBYg8T1fupS9aOaoxmIITXa+YBwRb7y1InZU5fptI2N4TNgLo
MOGswnFP8Xu9YRTWo+T/ApWQHeF08VrOUhG6qjPKJFIbUn3YdMMMh2JE9uG5pYofMsh73ai2DGqs
jYwQsVnEihip7W76aSMwMzcATJGZ0AZn2d25vWLP5f7I5if8by7MxPq1veowe7W4fjjX/nLJSLD6
PomDQ3QMZl4lhfwbpS3jl9agtGq/KZ3tKfBWCnlpItFh+eTBa7wWBDG2M9bQHDtrcdzfU1Qfc9WK
4SnRlMOGlitmbTqJAJzn/iT0UuRpDWmGE9VLFw+YCxYPIlfSn+hz015h6HlmhsA/N30Zn8ukdf/q
lHk3cmCwuPGuIkPxLhAxg1LvWK/5ZUQFjEMKwB3YsfYp8TCt0tj2pUw6jQKxncYj4Z21TYFGoL7O
MoJfk0UONOsI1ZNNUycGOdt3FEp1URq1kVckPxCpt63oLrIBhvRbz8XXrZGFOyZvuGrlLAFu6+qa
Tu54zkEP9CEDnA+cXghIkr6Sh5lw9mRx1wXJ4tqUygjW5EtWHYELuofQoLvgUG+cTznkul7ImxTC
0SqFbRpw82eTPBb2VtBw+CXPslhQMZvhFzgZ3Ytxhwv4AlEDcZYMps9upEVgMu0le4JLgL4naATb
kxdZW0taRBjBWxg6WNHUCevqJbxWFY9sIArZpRASlGlFhTvInPezu2ptKdF+XhN6UHlwGCuSd5ip
X2h+jiaINfcIiVGCLBaMThd8j+RlH6OV/tmOF9axHc/0DOZBOtZguOUXSX5FUbPfuTOlAu07c1OB
rOe6zB0d/ttQmGV/jGK1T5s+r3ENA6ImHD1qWcPEX0KVjdQtu9jOtqC1xkmZ4+LmjMsuZVzQ+wdg
vUzXvJARxQuGTjqBZYFuw/dFAef3tNSQs/bD5N+mQRfc2N0NBD8ezFsI2hDPAzmEdvFQBUyvAySn
3lZlZnadV8Eo4ItPSnOVGR3ApXIvBOAqlpiu9olDkRvb8pEfkj+BYTCygzOmgFHRGHCK5LWIqnxG
ZSOiSrBWoIuqMPG0s2GSsjwou48jcvMLLP0u7IOda9kjVHNJ4ryhU04Hwn0nghYwvgnRm8FUTJbz
FvlvADRpRgZaqzgJYMfyf2UxroiQBgq3wAO6u0MMrcC8f/UrZtsiJ1behAtDIzimSlM3kvtrfBVl
bj1YYSroNe/2eePpbmhlDIIDkVX6KajcexRc2VMkJTMcHPCRSd/vghZJZpKH4a9zmSNfAhqwKQby
ytoKwqe1JyFmVeP0aerSF8H0t4rGLs1WZN6RluUoCvdZoKQfQ1ZYU/w/pV2qbT4XJWTEvuN0Vkvz
tMrb63Qmbrrlx0CNo3AVxCUTQg+eG2u7NevNF9LHHMVI+3m+GXbol6KHQcFDl7IhyQbhIbQ55TZ8
6dzn8/kv/oIlFVCQ8RcyGzdlw7Spw3MPG1XMyYNJ9yB+HgVAWtVdDfJTWpm1ziXcQbqSA1wLGuD0
CoN8OhNcLo+bJPUVb0uFIPcm2gQPwqMIYtXitx4L402mM0V0IBUM89y1kT8D2eQb3vsqKdX6ne/P
GvK/4RC9xL1prjDB8bQY3jj/B4TM310d9nG+grLXiYAIxviONS+YdIH4rfz2bwHmCSg3DfJcMLmk
AcofDE0g9XZHQDPc7Ke/f2GBQezltWWBZhBQP26RkkHCpczKnOznYC0UdaTRjn4kPDxPp2umJ00d
W/+9Voi3uxrEyVZh8QmI8KvexSH+NYg8NKwW95pA8C7ipXA7YYu/TlxHCcpUemrU6JAazynzoPQh
8k1MWnsrt/MFviHX2SWHeEgS5YcfSsG3SmPdtHF4uPxTXFGktQwpAo8RLPgwl918mwwD8j0jCpST
Vm2Z3iCvVEutPkc8ei+ZQf6uu85bf5Rw4J+RHnyFQDi83I6LZlApM/S7ySQhDZ7s41u9G44XQ4VH
CkO3iX06FbjcW9Y04ReEspx5NJ4VYiqG8u+8RtQjQhdgfgqk8qYOsq3fJCe1Gk/x0LnmVyQoBa3b
w+fTg75vFWrD+3BnwcwxbmdfqYwsEX13kXTRew0iGt2XILUG+C8iXZwjRrUc4EpACwqbyY5PgH34
J5ilPp3IWAmU3kwUaCD19+17+aTFLUdsHhRce2fpgguzvt+iuCPop61kK4+JTsrNZh1SUF//6fjE
4+B/bxFFSnLEgQG2ccwkrPJFtLSNZN/fkqDS95q4aqqpIAxFpgbkr2VbLBkYMnfNER79X27y/f3t
XzWQYpBc7xokXkbF1ZPM638RCFqay/ybMdsSGBYIJn17EW5kBYJxaE73WMepZKEWicGb2eQyi/qc
JnqDSxuCsxGY4qy64LO2s4s5L67QxKDSsKEnXqv8rGLf04ay3f4pYs9RnT+36FUAyLdw07ggwI3f
KADE1a5ZOCO7tyOn2t1VLm8LgcZshxFXB2q00aT6YoSGvQlR9duynnFhAXnvDml1vduGYRK7thiT
AueHn5yZGP6YVgrURxcewLQI4juGyWCuFXSKL3T7SFyg8iL2lBIIRg88JsOvkoP98kwU463+0YfZ
+e3Ijv7Lywv1Hkgwd5JDUmfZc29E6MjW5No7bwsQF43xgJX+WtQvIyD8cVDi2w/kHtX3+6yomQb1
Z2g2U4qm87d4xovo0KC9d4A+wiibfYtOrvjiluz4FWr3TotOZvfeLYalVlwi/plyQrOTpWzAlq1i
/1uMivzyKrMJ72HjGphSifxHnjjbKmirVPppbNsCg9sJodyQCNrKySiAcB6sokBforv/xbJknB19
LlkykSISMLT/UomptdVqSiQGZs/ZxcylyVqCid6/nQMj3kLDUV4ScKfczz9V2VxLVKN8c6bT7IVe
xJDCDgjrCEX5Awt+4so/u1R8zoP4tbglLhpP7sFI6aiMPXpK31yuCAjMhZMY2GyCnPz7+RCszK8V
zfoijj34dLLkk+hbEJ9lLhIuhYYI8pYzMrZWgVHio2Vu9DDgH9IJQVSra1MTcTsZ2/mljJ46gGmJ
sAq3cUHG0FBmoY1GnX6WYUr+kBHQM1n9zbYJ4EYOnmwHajQg9/CzpoMNPtnj9CVNAmlu8U2z0bus
kadVnFxxOUtm4YqPPOLROeQ94FW5J9lVx5h4+2KKGZd7Ot/UGR4fjIABO/pfAdDJtURGaJIDMySH
rXPNhQtFhhYeb/PfPbGWjs4OLjXJ3FHmnoswwuXws06A+QsAUkMhJxJUWcGevb3hMsPse1Mhmaij
aFxQkNgHAjdb4nY9Gb2YAwpmtkypVoVyPGSJ1ftC8VEc6E51mnxHrK3ZH4nb07wOLXKF/zefGwkJ
tOyOkBFgQvHMpzmWQu4MsRX9P0edLhAOAawQx8QglkgEL1bLTLSYPukT2cPHn276L+46xeO8tT8t
yJw133On4iTQVK9+hT1KzJJiKcdB8Oi9HSrHGmYZbu3uZswZXqXQa2c1toV7ptJn3yDQeCnp0GuO
/jbP1f++GuBLyspGgoIALTs6v5eZ3XLEbInHCeT3PuQ3KUBLDSNsirnXz0D/8aT8n/Q2/g/Gjxrj
ulcxMprFmGMcK3Iefjal22W9dr9PYzfCg5XBgUGOWIIbjx+lT44n3lVAvemOckVoFRAmS1rSnAIP
KXhejwwFynD64nh4W9Pr22fcESZMAQKV5q//wl494pX2NsdeJInD9I8O31/9fb9n0tDf5gi/VYUz
ixzlvpesOiKwsNab7pMgPxhADfK98JyBPvkkGn8QWOfw0LEBPMbf7ltERD41+uq76+Hl83u07LpF
0vgGQFSNrhw4I6QJYhQrSqTb+PE9wvdFVlAWZzltOgTB9YDtcmoCBOwWO+ppGSKq/euSD2yjGgss
c68mVqdyw2sfOZZxStiqN/dvWSsffoJI+7Kq3Hn4uTJ3zLhOia/qo8F2FZQSLJD5PuLQaV36pmfO
AMAx+wtEmeXCJPGAY9SEfYMJH6xCEVJPNfqWNjikuExoQiaqbuor+RDk0L5eDA8vRIkkN/N1ZZI0
TgLIceLDmEYG+7KK0uuxnn+F/RhbInW5H2y+bX7yEzgkZLsTGPjt6eJM2pizFgyCi7gwODAmlti8
a15T3X5lOiifv34AIxqZ/8AhImlN6+rw7b+/NS3wM0JjabP6myAYrFpoqhWx84c+4gO6YeNn7Fo/
8tCP2GO1/20qUd2V0QLNgLchi78DPKvOe+sJ/mbBGt4XKe0InXxYlOP+hC0wtKdx67muFUZyCgqh
N7onn/Ux3xCu2cKEL0CE/R/5DqFX25zYydn/a+4jpBxe7ciBeih75EkE7OrckFy348JdkYefvxm0
ZQ3BViyQvktOwzxPnpvt1pqbndksdymUYVb8WZaVnnoP4ehb3LVXawWc7mQ4jiie1HrAqpH3bLzh
eQIYFQxyv7vzxj9wbNkmEkuhgn2nlneHggCS5U6mFJMAWpkAQ0pwz/5uAV40jsaBZrX4BWfCH/3x
9dPO6hSwzP89Wazl/Y7qfiwO0UnzuI9oiB8XqBaamdPavurHuuFf7dG+XTGFBZLzoB0JlwgewDWe
+GYLghIUY7dh8JtUPEynUmw9qD5lNqZVjGj70zz9ZZuDhiW7VvXJZwDMYGY/8PKMk6K88RIG4f6c
TWj9qsXBtaCs9YRDK+11caGXv89sMsh0n8MVARnQ0TGH6bHV1tOJ5eqngxB3WsPkzWpqmC1++iDS
cyngUPOB7FXAyX9pBjf9VH+fkrXq153zCkb3st+2AtRGd4ugRfjaOcXQtOivBugC8mJVLIfsigcr
KvsLje3zjkxSe+3PDdqSry9IrAwSfM1v0/Yo6l+sUZt/hVfpMKoTAzBfdxSNHSHrCw6AGNhxeazj
KjVhtVY9Y916SPBNh3dCxP3zztrf+wJXFG4Cokaqp9pMxkQJb1R+tz/c6I333DJOHN+madxlJyo1
PFJ+t6RG9nFJp2Iad8tqqvG5zABHlxHOEFYTarU+S0cxnLjcjtHamAA+2BcWYsHJ/tz0L5b0nl9L
8u0RElYeUgkM0axt3pHOYMr4jM/pyMle1kw9JasqkryhHo5u+hDm0X1Q0JhWAQX4U7LvDQOqDZwa
XcVlkjju1nNvJTtMbVlUE8uGgh59Q/vFRhi4pplcl/5DDuivezufnONTsU/kk5cNahBgr6WsUSXT
+o3VW4vmK5QxQgM+OCHdgAjKpPOovbGNxqtnf1UPkkui6U8/TCSqP0vxehh4AJZ8NjFKr8dLfTl/
Bjsqquz1Oe06OiU3pDXYoAvCjYD9nbL1AZ7nzqNF5svnN3rKnOwya/PqkSGooRdjTsVwTfWsaFD9
9xWVgq6WvP+R8MemCeBquk39NLL0eQBz6A1Yt1H32lx0gQEAhxR/RWB1WwsFE94OxvEH1lNblrvz
JmPl5GOjLL7j9beZSEs7LWPigkWP7dUo7o/5rFRNdc9kGKoXN20HnNqxcm6qzhOUMKtRlHDMY5gB
LUI6i76x3m1/g0LeRePRFZ+guGGda5zpA7QDsoX1ggF6qA9CL8cnlNk8mET7VeWhEXpoU8vdhjWg
Sggfc82LmGM4FOxqqoJvuYRxltzUgjZTh84Mb9G4PKlb8+qpwpDVrqbleb9x3DL6GKjC4LMdSoUu
EstevhC1Ad0ijYjxwgdeJ+yJdONFSAx63Rn8whJiisii/zDRNW5h7tppzbi8YTE1gPZvIe3VA5K/
bV4NHJiDH6lcBKYRpcVx+bsoIKP5Hxb4eYLlMx9Ptr/Q8qlR1hj35Qcv2PP8gzSrj19FMvyKEyxQ
PcaTyXK3KDcUkVB5anPvYZ2Mvr13VIEc8DOrpG5H7R3aOMYW8pvndrrPFoxCPmCFV65hpYbUhSsO
NaFM0cRWf1dKDOUsPCSM3Nw8+QBHcp56+Zb5tuJqVAxU1vNfIGw+wVG/E6gyxzHWOoUpGXaBLStE
xBLW/VJGsNKF9Rc/W6DJeTDjS+qTz9ReGAZwxWsOfhJ+13zLDobkj7hCEOPr7QHShxbeJyW1NAtS
Np9oabBMrNPyUEr5pmxbKn+G97eqt1iisWG4WfM1k+ZsymZN6irtGS1qHguVC9lwsXXK51tPae+P
VJskk+wKV447BYyOBH9T9swWU0WCuJsCfdlaxlDqvXhXUKKB3oNFHBwbYR36p+9Yv5ySd/n4J2dE
bOYDzoYZbiV7aGzMp53BG7LdGasZ3ov/1gY/v25Alwinni2DADgyAy9JPup7fr2ULa3KMh4eVoGC
8GE9MM+455tfsJEjWx+JSrgb1nwhaUk7euvC8Uig1C4IlK39hAURSR79wzboKx033KQAg2Vdu2WA
k9RVjhGdlgidzKUAdQtMIoDSY4ysb78bnx+TuoKP2Q6Yi6/zkDphLJHN1TESDzj6sw05TumZMFKT
HcWcX+Kz7EU5hOZ49chHRaVVcJ97igRX1v4mp3PkFMm2Olkb3zWbeJRMe8J9g3/tCOVrDySWXieT
jct8/a3JoNDNyJyHEFF+In96a32mBV1o9U5BaBwiMKEi2S8xJroikiMmBB0S2RM5DlT7x5qt/Q46
MIRHdlLQckx6MWhQ71U4P6Arrmpz8U4gLKOfUL2uegGxz1G1jiX7UaxWbYGeCy5or67rlL0N3/N5
1HCB8tlLgxteEXpPSckIZYvACrxMCIx6hZYFXRVmUYWtccVQGu/JFfSsYJ0csRQkFI+ezp7npqdK
dCxZ9oneB14GzenVXBGpK3l4+UsTv7WaTZKlQPmmmUUC0+kijsQyE75FQJXz3zkHrI4uyt7uYIst
WMxyl9OhYtgWUdxitKSJvvtzz8q+2h9g98vWG7Cc25zakVBH57ppJJdeMFyq2A59IIPL+2hzYV03
MuTyO+UGMbJjSCCFuJ11Cwk0WGT3UNUxk0Dk0wmbSmKJQq7q+noM/i0z7jJGVEKkvEWSqYK9K/FJ
CLaDpJIrynh7EwOnJwEMyp7NF+b+fxJi0TJo5DJm+shqkN8ertu05frfOIi2EfqY4sW+m8XyzeA6
ln6HXvR4b5rTY59JwsrBqyxjVSP8gZK+1J3Lz2++zBbqWdUlbjATVnX/HA3zVhAqoseAygTu0Hph
42ZvxE0Mw68NldV0JJ9YzzVRwMY0nDAiNJ4stz6QoDBQ/Bxw/5mvWPIXKvNOEtpU33FB+MeyAGP5
Hx4rzCnYv6SAqtnCNubRimp/id2hzmIg8VlwYwKaeDOGL93L6w9ACKXUmwMzsrDLsH1xg3EicvLd
x8V6aQl+COolaudGiplTBRlKJbEYypr4V6z+OxkpaZQjaxTIHz7MPeo3rct1QdqitDBF4OKb8E9W
WzucQxc2VoOHaRsdge1KDlHihzwqulHfFDqFbDB7wwL7B8Ar44f6sJaeQc6Ik0HfK/UmlxVYU/pH
UVnXThPvjmK0ToSiNwZveBxzq0psmbhtbe8jUWMfTDvJp4m8yZi12GAIim7umcrRktk5Lhv62CpZ
9EB+k7QnPXus2L6Rc0uITdnd9qfLlv2c7A46SS4OAT44oP8rE43AvgNywyRheinTe6gVApDL5Pmh
vOe45ovWl5vJ0h5OPq28QyjLgJCYBToCC3H+VweFIJumYo0EC262SkcJBZGAUUTZkOKwlWi13ljf
j9sVKxLdMJFsEm+VoH167dyNzoUg/xNv3ZCy4mF/lETcry16msmdxo5Ewg1salULybz95B4sYRdR
4JkC9eIOgN9OMt795lHa5gQnUZ92YUOWfvEwpUIeXYHmwwQmnDaXrFQcNoYD+i0D/v4QnRU5BB4F
g3UVda1TisbF13rp7WpChpu8YhvrYTwuG/B3uoRL+IDbA9EoI3nBRDKWPnPevqi2ECdmYi4W3Kmb
H6CEZkh6yycMHUSLJJdYOHGdK9SYu/Dii2NX3eYIGghdhHxDTFeHnp//XCwNWrJuXFplZG+XCORH
VnrIyFyNNXOkESO5m7GyasR8qK8BF1K+QF3vN2KBbdTDglz3hw3VxuFC0I0TBExfRKaUj+XTw/9W
P1vCo89GU+nLPcALJ7UDLzkFgSsqpWsX6q7bKUNXfOtdQ9iJxL87DuM1Fkmr75HQTWE+GI2onyyY
PVEziATE7997jtswxn8m4/5GV5CW1abHCWisuH4WvGlQoGskyvjX9PGAahSUYhSQ9EnjtvnPUfpy
jxK9hcq2vGXahVtRykhqLGmTfJBjRDX0SMP1AFaZZh9bhNEvbWxQXzuz0+zu3zJvpme5DDmM8oKt
/kxE9Tr8ye0g5mzHpkCQD9bC1+mq+qFisG7emXp0VB3YOAG5wZ0EUaeiFbyqOHrj2+LNrFn8Aul/
WTbZ8XaM/4jppIvENsPFRDRu88f0mO55vbdEfSD+a1QJtS1T425uMMtqHTUmTOIuy8q3zugP4fhO
Ltv7gcpZffwvijaOU1LnZBG4h3aiZnfOf30Rb7z40AhutvvEwdg0qJ9PZAMfofcgsENgPNECGH/h
ME4BSj+sj39IYn54EF9VmvXV4CUvb0WoMUKbjOms1Q3ALqiF2XHGvjYOlUovNxPCEOScXibtEmRf
wqAU6HwuEVw09DuLEdWSR01NrOgSq2LfvF9CYZWAw1SArrVkpGn/Q/QlsrOet9uTjwq/hE3wpHWN
+viW53NF82zRey7YW/LmF9poZY3pqkAd/NQ8MKOdpou1G70v7CDbZnJLDip94OmhLtFV3thck9qx
yovkNdPBkYdPL7adpee0saXeRDswgT8K/opv0SgmjLrB1JxnFYImBXbb2WnfanRcomJLDlJimyJB
4NrUXecWFlKTIHkycLRM7hWgmPbNBKMNuzjFgPR+7XtIVrAKd1nJ3Y1w+zf2eWDlH4XkFuItJcyn
2h8Nb+NOlCWBHC0Wpzirx8NEztU++RSkQtaI71tzd9fB9pWcn5Jb6KS/teOWB3dn8kOwfszDuE/q
uhoTKaJW6yTa/kGsW62+zioVxlgdgfxXPWqQrCm9bNKSS3FwTaaOQ6ijrQ2Y3kgk0YAHK+X64Qos
g6x0FZYS7qrpu88SpsnttuY0/7WDZpK3SJh4IaLc+AOz+1czMkIhGJUc7apJ95Unp0Pzh83LNBTL
X/xI+I4idW4VbZlTtbcxeO6MPv62UDOlKPGgujq1k8YpLmVGLo1VVpoEoHP4x7qk/VKahO4B3Uwh
sZ2l4HWJpM0ki5WadZaM9gecxmQB7MdQbMwuwTcXhQpbzHYHgCUM+PsH2ZmgAquHyAudpot8vj+j
SEXdcSGaDjtRam5Udzyy93cLJn9hYeKynbtqUpLQdvIS4v8O58ALVl8sjuxuRuqmEfDQrQvNR0BL
ZR2vdE92/HZ8dNBUTL6lfjLgOYofVWxRWz/sfvLEk5Pntmj/fP7gym7uYRrG2sERc1uDTrEBrVAt
4E8qHE+Zg3YfffyAPI8Rjey9uP4DVSLRdJw+OjltQE6AxZquqNZN95OID2BTNCCARgQy8uReyaOL
EW790dejprLtJGW63eqhmPq8kI41OPrAnIbewSysBnXlIEd09dVi7MFIdyfmy49ufeaJ3MRu/hMa
2cvR9TskfhyPHGlTkP9vT5i7C9fZoziO1//LpQC6u6A9nN09s8MIQuS9vbdWAIofxiVEQH3eFTMI
BrQOEoKqIU1XIrfFpifmme0q0hlfwdRhVYoB7GdjTwd3nu/7KGKLMBKKYUiTGUoO6jqo2+L/Bg7V
Uhqx1vwgbqOGM7i4gtuZUsLHhick7k+rfemd4XInOAmAiSeO3rcWn1Q/R1vgDM0Z7jB/pehWAzqQ
JLnMX7qW/RjvyFF3RpQHpnzfh5lFKBU7sQOXlX+hotuuxzk3V9eEicaPX5FyZUhfzrauEw4GdOyj
m45g+yNAMhOR6jiBhsQMODjSzpDy28hNGeiO3qqBjUXWOYmtJc28xtpMiQ8YCV+et+5f2UxtfVZS
McPEQZBJ/Rtz+aId+o2Cr2HKSusiIEPkY2aJgvokSWksj6Vj4S+QyCCTphdV1jRCcSGtHtjAFaqz
9r+6GB6VUftQR0rlwizhN4Tb19o5PtshlCDgCSnI+Mhe+FRBZxiEfAzQzSb3k5MJA8QdO1a6iQrE
C3vqM9kZG9NE+Z8SIvMjGEGamoTrBA2AGz/i1412BQyW9YlYWCaZhVmK/dV3FySD4bgZycS+znNc
E7svJ4CQjydKhwtpfwrAEMDBCHJaUkZAfH7eQotTPhcbg21LXBGbMY2myFgH1w+HASbRac6KiN1v
z5r557RuYAS7JxtSq3n7aP5UMNQBeJ78fX/jyEhVb1I9pqcHpkT0eBKoNiWClZRnhNyi/lDyewbu
Qu/J6+CCg6usc+P+LTMuVVzZpvFRTP/oaQ7uMs3APxqpxHWEnFanUzGCFAQWpNn15wOIiza+Vg0S
3YumGjVI9dlwj+39mXp6FhtELtmE0Op8OcN7TXOTxyCPXjtVgM6F3J+yhftWiWGrOmQX3+OS3hSY
zCIOxZtIbjlyF8zP9byys5Z9hRITRQJNbDyhnA2taVWKY1cLmZZ5QeeG4ihYotTKrCdD9trMJT2j
HsHIE7Mv0W7AwyhZY7nX9q0TESTJzuUyLu0SZKWHNDHAPGdaxV9uC6hWxUwm76dYYHcOeaTzLroQ
s064HU+LIx52vVYYRn53vIKqjH4YLX/eOUh/flID9jzLxwecVuczSmxaWNU09q8lUaaoEYx4/Uo7
4KUKVwKc/LRCcu9YQPdcSg/248U3m38sAsjBES51g7ts0VAcEd+VysNBql4Ud9GkQxcLucIyJIYG
qVS6G5teR1BfCi/VY/JXLM/v80km6yFDTVsloxUpxvmbx2c22b/B0DwUHHcasMde0vEF9kZATC4e
/NQ28xK95/JQCYLHURR35y3NqOK2Zij+ySac8cXG8G3eUmcUlzZi8ZyVXwXfHh9H+0mBbZSCsohf
qJusILYadQ5+zmGXefn1b/IdDu3JVrJqt2HA01qa0QOaTH/dbFLeS1/RpJV4qfcCsKoOhktqqbO6
OVErFBDmB+nRzZSqwB+mNg2wgNngmzlKcNZ0FvydreZyJIBMUpFoy+W5Z3cRIub9X14iZ0BLR2Ue
QWVKTzqewjkALXDXX4CNwfHIGaw5yp4foTPZxvcldVcp3Yv/DeYPhDEozm002idjW9hN3soQtQtD
7rnuwhH5T9oSASereX6nqgVLpMHicECciu0i7WfPCaykKsxVR7PVvgAqan5lSxaiSankdELqg4ER
uA5R/zqnc/0XYRt4KbIbraWyq541Hni22BqBQlXtCBTw/0axF998JOaT74fIy3M6PeE718/NnZ5b
YN+dXk+T3ErrxnXsFQZPTVPyofA0ItFcvckmMco41OgMCStU9Dx5duV+Ocwe8wqZp5drWxJcnObj
2r2ISC6QQc7bkaVnlW9xYMkqxzXTNIXhIjvZlBhS18JtH+zIHAQEeMhHlp8NxicLeuAL/LnVOgzD
O9mLC8EATIXkfeLB8+XKlyJJeno5ZgpKIdV0173zYNNkzqb76qtgkZcqbjN6PIvzkpix5NfJlFuE
B8kznnruyghvHva9iH5DKitZjnUNjwH9fIzXrD7KaNqqtfXNGhYUR1idtuJu1sUSKcgPLhuo0KoN
gtb3oRrONqX8x8Me+eFpje0cOccaur3W20cPG/f47FXFd60SI4eJvty+ZxJFXQSztxpjOQ0ojK9g
gUY1SLP/E1C1qVr/U2DRZ+WVsxmBb3LoyWaL1r6A2OqtXKwF3aRNZPJeoZtdtYdsso0mLsfYHzyM
Im1YB05N5VeUKVdTf3A0r7bBQJ9hJmO3IhXyHc9SxUTnZ/m8deOWrAjjd/WiRSIg2llj95f3U8Oe
NlhVVwlj8KOq3NcMuKRjVhcwSyctdXPQQSEerM4F6g0abfs5A+Nk8mpM3qfj5kZ9Rr3eG38uDoxq
ilGUI1GgRjLmbN40WB6od6CgWTyncHDPGwc1BwEIbkgQkXRNyOMdb64ohHHmdI3vnDZGqYdlytoe
S0Oo5T7XHLnY6a+QrFaPRgOfMKb+3rbEfqL9P+C/QpMsLpbpU4YcgWUU8yS4AazZrpAv+mFqXVso
0W/yMy//81rq+C0c6tcXlxQpUMm7Ke4MlNDHh3cOdgIQpYkPmPRJVBJHsCsYnvFW3DIQgIJHLwKY
Mtz1zqyVf+BjRrXOEE6aZEoLUWUFgSmAhglYq9OO2uFVxokZDRgAuUL8uEXmPnbM+N4tV6alBZAj
NkXkAwlANBiSFB+pehk61a7eKm58xp7bbzq08TsbFBH5BIKiZntnXR8S2cDZWRuR7595GtIrNeY3
1kyj1NgIl6lprciIAhFOtiVDUcp39y7tcqn1NFjzOJ3rN5Naz+xqbXgQxGkDElzodv+RJ/TU3xH3
2au3DgATZefP6q/w32/vjjyCFD7PvGsQDmLkmdP+Jl8t7uWVCBw2yypQGcrmPtn9V6m9eFG51ZJv
7C7UkH0+rjSc3SuWYRHVIv+wdzQH58FktM5UMbG9k2AZGoVtHX+kwZI7eIJDiAUesr9M5xfpuB40
Ii4MrqcWEK2gK8WUJ16H5ab3vehaodUKVsSXX2hHUg8XfJiZxksA4KsGrnYc52OO12FGzLMVibT6
3yaSmF6K9etd93p6hgUxCeWWiRXOyvh3fvI2ZJR39s6GelJ+YveIqIHydJa0felkwgWUh9o2OSwN
tnKrPNknclLb2/wDfVJIRFDvz6myUqGwBu5+y22aHsJ7iESmYIcPGTAzG7dHAdLkX/T82/mA6idy
7FvmampuozWE8GCTf8bmJdeyp+NI7riHMYocCV86VhfGFa783KCqQZ5yfxupvdAWl/lWA2HioZh3
j+9LQwx0/GYr59INrgKdUTJmbv9x5PFSbYfJDiJ4D4YFgOBc5FgwoGUi8jkmmejjm/7x8P5IGAu9
o7iMBx8eVltqDBvgeQw7TXVnjRzAcjh1/LX2uWJKVnxqazoLUCqiH5lGbMEHYTCRVXZ724qmAAfi
ipbQKiM5CXqSePJwTH6aGV53uLGSnoapEiDXWtLhIJ41MazR6Xq9cU6nrXvq+S8nKP9kVEPohmBd
X2AnKWgp88PiOKx/iL6oy0wKt2gPQlwcdkgX2X6HgWurfy22UWj1azFCPpOjyBmxOV7ypQ1DFFcE
shANUYbz18inLHy+/gXBPUjMh212MDf+HVNe5sIGVzjHAg0RXlKqAQ5jvaFQXcgylxEgcxANlsiI
A4vneyVT1F096rCqaUPndZWDHzZPgqPix1C3iikmv0sflCGnHHneiYuMr4qxK81p891yBYYv9Nv6
dmhX+a4ulsTXUR+qK5LxS9pBp0ycltolFiQp4pR2lUUxFZXxCVD4UiEhCch801u5/8isXFdufefC
e93nSKXdioRBs1R931fs8XImZ1Nesd64pgacyNRSWpkHLUXUp5dM+30OA1HSpAewtKHyoYvy95XR
BZ9Ewr72zrbBIYhtlYSN+l7R7uyIUIHM84wUvV3XFAUxBvnMs114L2eqmGn18jy5JRA1Aw5S93bO
WKPqv+YTUHXSb7+CHtc/4HZq+nKSPJwZPxm1YoQSSJtKq5O2vRM/qNSFDrrY4QXb4tWBSlp3mprz
20dgLa8TLOH7XOsWd6BM6jbBC/zZLQBpVlBnjnMoWB12BCSbrTTEH9QNh/5G2KE7FsiWwlTvIDhl
8YnNesufYsx9ClS836m0w6C/h3fWgi/EZIoz53vJ+S2EZWgGhpDd27juPJDhisSst8Nzt5q91SPF
GYdIbpUsZRkHGlgg+L6ejGlZhouqlEDl65WUQUw3F6QMV9bf5mAjMPK+dqDv0e1tTKRCZkcscOFH
8SofvV/Y55osrHkBJL1IPNrMUQkYvyLGIaimal0UJInyzGc2Qcf30CoteI85eQ0SO3Uc0uqnGCJa
zP8imWmSQPQvfctmfZncJeUYiGKJTd94uNWVWIgGGUcjLlKxxrxUE9A5NLZ4PkPg9Ya+WDtcR1S9
QJDmFvgknFUuG7eNrkgpssTj/oeq1vTjAU9ljnMK9YdtfXslUl9OiAp5aOSKkBuoHAPF4n1Tp0fx
AVufSsBs/xKeifEjGLDR8QeJxhSQbb9mmjIZp0ZawEeJ+HRXF2Gfh2aO77PcaQHm78pucNiEmDbp
yw2TjeB745H3wELCUp86m9sXV8HFT/f6ngNVZrCVX7KCJ+8mbhx8DeamVKDnXqbrwxvQtGHlQJnn
x5GtqC/wcI4FgoYZv6rec1fcdkUYzK30DdSZuu3KsP64dzB8/CggIW8++pQOAw97Rxng8o16qCki
lkxsCEpVW6XXDOF8bTjYyfeGGhHyTc+7L44KMCa9bZzfNZZDxnEVbWiOcUlSM6qNwIrRv6SpSFIf
Fk0tdgTic1p2XsNMTLVtNOj2soqS2D6j1W6uv7VvLrB4nPnKTImVfAZFg+FfestwPE6fuo4Xzp9B
mCNbjnBkcnVD2QqsvnYdzJ+m89s45i7bwIfs6/nSWfbE8nnGNozrACcO6tGTltSb4n1bNG/5eSl6
wHCj8Uizi717sAqgmavfHNwCy9hqmFoqJOJVlXkGO+xiZWgvHxcSk1hdOAoRYmVUdRIxgHOmQg6+
DcLhD9YfYRTTGf0aQ14fnUzwNUC62CH2w31jJ7np6Z2twFJLPNLL4sXCZCSqYSeF5e5N8KUhjWsB
2OOKGnwjyirCL7NN6Bla2J/nBUmMFbbuVu3ky8/uVSC/hdYb9uIzT+9insy7+eZ/2+FJjDJ1Q0lZ
b0eEbYX20SpeHuGhgxoqVdItdJ4jT51wVd6Gv6gCVrAD+7xxEI5SC5mxWq8RQ3VuVJLjw1I2h+oG
sE+ImjUkFeS/MiSzGxNmRhxif+WaeNqcOtzoAH5Itosj0YGnY6H+PHIoJWdLs5AHNK+5y3BloSDT
Knkg9SUJLTbPwJsRQmvLPM27RIf5rOU7QI+vZX+PDWh8tlPIACv4LnFxHxXZvSWfTmggihyQQfMW
HAhBmnGe4sCH83n5LNPtVR1mZnUD2OMDEwIoYVzhH+BMCy5b8tnrOjJU6k7GoNNVbJ+kO5xzdfLG
EouU8sMqHFZ0YuSdeNiyebOkyagDi4EhN+UbkATRHTtf2v8Cd/xOSfkeWGtel5ctsiQWlWfUWa3W
9J/l/n1M8czTwlcio18k099/lUyAujY7bFuZB2YQIND91Ox0Ev2nzUD9HxpJFs1zgBlk9SZ3JSkK
caZ1YpFtHrU14Fk03RQw1ef4hm/2Vnk96CGvjJ4YVpBJHyulN33IZpMmmTpoiIMZeMIC0jqkfMZh
0+2+gFwQ5xXgbgJluum0d50r80hN1E2y+QLhZZLz+vHXmUp6OsnqooWhc2JMIysaXU0S7VTZsdT1
S+XlqAPAH3GZ8jeKxhBXsvbhrigD63TCY8Uhk9qg+pwPOQUTs1bMBMElbidscwSfcG09DbpJneXt
66h+GT+4oV3ihxa6kmAmu7q2OAOwGonpn4D865G4a1YZ3VqAdkIXkZPHAgvk9gfZPSWYWuE3PgqH
ZWzvp3gfjaPQAEBvfB3hyvW4TplzuUJGpTKqF03QO+NZTtb7F+s7/Ss+az0ARYrk9FLykNpqsAIZ
7PDyrpRlLUcaWnUKJPeuZyeYkp2+P5tEUBIUtBb3A6fTD/TMUyhSHr+ATMJ/mUlDOdyoSNQb68EY
yF33r0U4es3UIDSlJIAjceA6bz1umwYw93YLaoMVGXldm/IN6RClwGrRXMgeEnFvmDVM/WTxB2SA
YS/GNg11Vm9y4bE2UwNincEJCxOSKAMn143kDG0AONZBkvg8VNGpsg3Ewesaj75H8FsXPHpJnp10
UX0iAEQmeV0rK5Nl9vLd+RS6YsKkF4IwNVSg5emhJ9qE8hPh4Amz98YPH2RXZPJ6F52A6GeEK77o
IjcU+Zp+agDLj2NFEaXJD5LZmDKOjnsB6g7LOvqAdbl13NIAAlOEdrh/nbMN7aynteEZl2VfcJUp
P8qc2MOTzFXuCg48Lhy9DdDpnJtDHcU2mCD9tR0fAu5uGZm9jysSDCAoKXlXnwLoPgLVusQc+w8Y
mx1tpYO17oqvK/oj3voRPURrDP61w3JX1Am+dVEpaFLZFQC8EKHay61nvjOqJhpD7jVwwYHyDvxM
7qPwrRVGCnx6jgivVoy0oisKSD+GAMHd4/7i87hlTWKclYbBse4u63XDtteH/fgHG9zcguL8Vy2E
CBHVeQ/WSyCTViYgNR5lgpu4BuHxNdzWfP7jiVXVcUG1xoIdojwcTVbNOcwMCfaTvIHENOpmYgh3
djFc2Vv89+NGH5Z8q/E2FQClGRMN1NJDBJGTB/zeJHdCcLAAD/V2S2k7mC52kPcD31P4YnDXtnNP
/w1INJaZ2uNFpr0+qBBxM9pOPLhT6VY2sJgVDdPxy0lyOydaPFn0lejNMBkCAa2chlsWOYL4vRq1
Kv+EhV4WydbBJYX/nH81FNmNgUmwiue4pbplPbZhY7UCnyaPCGYPgmTpfT5QfBvLuhktZT8URgZG
3tQFEUScQnygAvZTutgoG7jHvRZDpx9/DEgpFofNj8rwLP7gKxzIESa+QHERqtqY++VkfnyiCVla
nWIcjbLjzTog+pobSOXrc5kfMVeHk3r5hD/RJb+FU9HGzgzgYVTObjNj9ojxyGyhZkjbJSOHWURg
y6RpwUxN4YVAkPFsEnT+TNHocK6UElgCHERZ0ykAbSjmsZVmoNfRjCXvg0F9ktHgVO8SMuSbe4jX
jF7aSvW3l7jRNoTMymKZRwI+TKAOiM8N8kkK/h3CLCzmUGgIZnb7sMaAqi+/aNyDQurOkVxaSidm
OnKa44zzS0OmgzkzoI6jOV6in4ocnQuFXIR6+1zspbzNQxv1tCnwovO2APu18cATDwZAtvpPxba2
MdtePW/jmduoivpIXHggo2qcieUbg5gUAQ5JoXsqujWU+hNbGqqF8MsxEJBxyiEXyimEr8rIHHnp
dmhO0fGJD++6Zbn/9MfmsnYHMvUc1/P22rePHDIeXWqu5XPLTMSWuF7ftxOxW7/tzfM5jDIMKbX/
j9G27cdH//f1PEGW7h2ThmOHmYeYibM373/w8kBVCutOXm1dSg1HHrthe4J24jmP6W+EPnyPHQuq
Ha3CgzqhfgcHx9mtmna/Yt5ArQMj0SEDPRSFUX4NNjNo2pBvf75GqS3isqDEH4pOvHPp50EqvFu/
ngO14wRW3TKaYYrwrhnzr0e0v3r8rc5rTpEtBW+/8JPlbcsokYj4tQmfXUhM/HSBoD00GBcAV9dK
YZ3R6ZWlSO7XDCom7YhtrDZjNhDZ39qB2taMAyRej51n7vcmn6goGiWpLQDMXUnHD9hhTPYg8G2P
1oGU+bR7KUo9pl4VYX0OZ3n2m/otrl0hIsitiU/cMFOS3A2NOXoi9X2im7psSwczrgfcw8n5txqw
/aWfMx26AKbaY2snM2ryiCSN4y/d9TjnNZXUHXBZul2ihc8g4rESsgi0Gg8WUAlq0S7ggjWs3uGK
OZf/c62czPdiNlv8Ej+Jo/l/0vqsEBgIyeJJhH2+dxmGZLMq+dEjLznpMg2FtO/hFqgpozpjvTeN
5KcpnKks6rNTcaxUrD4FUo1vszz1Seyn192f/RzAfEz+5o4fwMRgIi6c+y50hH9znj/NetTAExJp
iM/rx5+bQlQHURbPQ/GMFxFBHVPi9sR+C25wxhSp6ORpfw6v7UQ3vpyYcgdNoYty6U72OSAkheOT
ABIwoxzybIllGab+MgthljMfigTvbD84By2ktec4hT2cc/9iX1hjRbPzY0zSb4ttWwNBxyxNt8AN
CCYxH3+Nr5C/UpQQluROsUk82HVi6t/ZVyejHmVeOrO7ESvOrdikaAn7yYPwxqZgCugfo0AXXa7q
4avQP/vbiNe4CWepEJ43H1bvS3DTUTih7i91wrO513oNtI+Bi+fOD5SF9WajjRm+U1OXYafLRjSj
QAZDbJj1mfZ2cCAhbuHU+Y2l94FMunf9hA0bLFdIT5sspVcnnJfZxxVPXrLphtweuwlo1GIYlfCM
BARx85GfOcd4bGPcA+uWg3t9gHtAQKo9dHkcJGQGSuuXInk+N6F2MWotz4WSt7t046osljRPw6UB
utEBwGOMlQ2iGCHqB55WtTCJLw9aZYTSYgGSg9C052aVRFph4+uyRAXnjUPkCJVMFZnJsMkuBZmU
dhriV5zB3kMlyT6K+cnsxOAxWR1Eh84F/Car/uL52p+L95CoqOjZgIz4yYLYWmloPSZL0pjnOd6E
S4UvpP1xph7LYxfF4MpB3BSNgwW5AZKs+tPKVw9Ns/8whcK/tyiHT/HAufIKMJozjYgrRNh83oW6
b/UJ9097DHwdkfVS+qjQITURMsMNdK8P5JGNcN6sHlrwNu4B9ok1GHJ6egJ+TwliRGbnH3I4QH+7
TxH3cm4EemHegZVaWUzEanypuFn4r9GmGQeb9TGRwwkrB2RdG8pq2O3zJQXJfl/ocVpiE1745IbI
dkifpzzHgoUWHhoNUCixN86heVNu1HvldbPxTNQ18s7Gb+tBXESh3/enrYYmziadLXTdRob1OKsZ
3Bv74NqRgOVqJDROcEOjIYqM5sPf0k445KCyFsZdQlgyDwy9qDx0Um5yHgMZ2LMfbJly0hsJ1mAv
PZiEgRS7CG6vgyjXQlpE33nCC8GIqooQhhai1oRlAfIvPYRhx21rdQkvbpOU8gY0V349ETsTQ531
iUHf3VdDi0cjNPNI8Ulp2yhNsOW403Yjh8LqVEy1JIKy6tucZR6U/8FgrMLsbXSukPSb6lkTQtpb
62FOiL0ciW4CiSW8ONajmAkBLrLWwLLNdRfYZEYj5cKTNX1wxLdOxy9lOxQufQYYcMkhCOiv0Pkt
eTTJRQGTE09iRMoGUiAEJ1jJb8f8di3bIcdCLEFCn5+NujHnvIQFlp1D08dM2pLlyCfJOSSzHHDf
F8Q8GYpVSeNu1oPhryC/eH+eEoUhrxiWG1+vcka0+glMOiEfTqAQ/z9JkVSpq6aCNfHDyZ0osEri
Nk683ng62QGfsgc/lNUfLRpVSdsme3kOvGFWhfaIaFYVdZ098sQtTcSj0Lgnji22bLbwaAHV6Gfw
hPI1gE8QiaH8ucr2OrVx/ADFfQInqbvZ8xkyOwIyhX3qx8HNDFH1u0f16uZCwN2DpkK4CggwSBWf
CWcpcptKYFJlB9XPHPUWMax3TRcrF2wJVQRHaWkrpSP4XxTs/RDftZIusZcg0NVC+xvWVYdO8TrP
Xr3BYTmS/d8Q/1E2lxf1p9Aq3wmpd6lKJU+6N9s3gjmvMoUdsVaq8txLi1F1A/lnvQTHSkzPHw5Z
EbM9+LVQKG/RvQulLGzkhipG5tGb+6fQPHlq7xPSDxk41K9NmGHOph9Ufkd6Bih7iBG/duxmJ2OF
aOfk5MmmPFokJj0Yn20g8G8oi//erU4GY23L3EgVNs1rOn3iZj77TNW9bcC1aTmIPOLLMgtRUy4H
X5YDQeWqzaGFPkgxbxi3AoPCDCPopoe9tecu4na52D8hVVpIFCkBC5U/hp1tK2HyonOmX1EWxScL
E9cyOnyTZMOFTt7eFPMt+kHBTS2c7G4Wcfo5w52Y7YZLOwuWML8XejBQzI22y06MlUbkv9fzxIxy
vlmNmFGjGf1h77thl2dwkgiDG55u5djhVK0/FYq/o45bRH8YMDhBocIlokaz/TbUm/C2z+Jb95xR
pjREj34ekt9gSo2W/kf8CQSq5XsfI1mh0yI1w8DhdcU0eolg9w5YcLs9AlrLgGmd4vS5X9myFTGs
L2mvK58RzaAtHnucg7r13WbhwVCis2Wluv4Neezq1dWvuTdUyLWLr94RBIuOjpE1LVATmMii42k4
2kK51I4D6XCz+MuKWUAXc7xFP2v5OmbWpCIyE5ok6Mz5L6nGzrVJvI0kOvWOCnpSLUPe7HFFca7O
v+HalDpjgBw4ozYuEvBT6q9C/7n4GPfrvYxjlzy0Si5EdwfwyPhsbcN2XPq/ymYOiJaQLnQ+/CAd
A2nHAja5n+lIcpT2giIE4AiBvN9U7KW2qzDjoymQasGcAsXKL/DKDO/Z5+U7EGeWVXFAeh1W4LgW
rWZX5yQytHnXFwZz/x2CQVsBLOVEF1jj5riN2GV22RtUpeie8dGCalzZha4L2GmnvSvsNVfZHUZ+
oml33I4G2Pr7AOEo/IYyutqPM+GcvVxNzmRaQMtyL7ZTskCjJEZZhXOmc22xDt4tsTYuCqErZ0Y2
oVjSdBngPrrai3VheJRLHdCRHRrQd8oKJ1oy+pp7olYakIL/Q+i9577k1z3sapHEj9m5yPiNBsuQ
87SjsAAmWzE9f1ky9whVCU/+GrNTgjPGwpvoRsJHSnJcMa5dVGQ5BIgxyFKF/U1yaSR5ztaMoPah
2zXUvqceaEJW+GvP+myh7k+mbgYoc6Xv11Bcz/dV7lf9OgPr6V10dwuRn9w1yR9p3yoxhNCtQwIH
gXCSahoHT9fLtw8L/50Ap7913j3su3Byd+mb/h+oNJ5IOZ2wGEgn0kaR83o9Oo4Wk8MFf2mkCQmW
1qQ0EJrQAl3jT435Dt/6ZaUt3GDdMlAXDmOev9TxZ2UNgs/zlPIp+HWj4q2pv/ntFPzpDA88xfky
h4x0mcL8Rbf/jU1+syrIsJl2qKpeUPE+VarjSQzUdff9MkxCx0A3UB6FKKjFdw05ydYww602MF18
KWWK8fisxi8Z826xOY3Bje1qX0/ieBNjJkAh7n90hYq/zeNk9lF2+xYroptqmgk8MToForfsmJrQ
VyfeGjU/CledTdCH9sGsmqnFNdPJW84IjDAdAVjju2bP24os/KQPLxGp5SKpSo/VeKfR3FYEC+BY
g5M6TMpLsgNC3EsVQ08SwiKEFq3i+DThDm99TBLopBD3TttpKQaw1W0oiMPMwVFz6IP4BGWDHdj6
IXSHGJf/Vb4Z+4T8dGaGJQECqKN3xia+oXcyM4OSnvZfLTP/GLLVdSIMh1NSxhjWh8dE2Gfhicaf
PSlWceTkZFpnnORwrwXQYiI/24PpyqWvjFjMDH6dQhOHXlSIwpvn7XhVhKB1B8rIWQVpRT9Z8GTU
fJtCJXMCbuN+zRzmn/OzzQVv1RKVgSMYdIztmWAYnBITR1Us9jL5JdMdmDaFERq2pg743X3pT1LE
PawB1P8hn3GBsKaSidlWK4tCRoSpSp5XTxvjf+sxyM+ap4M5bQ9ORclKClT7/i474G9ko0N9/7pA
XDznqjVMvhJlDlUFXLxB7e1ipqpbBBDClmRdvDOIuonqlb7bRn51T+VtgS2JUEIYlFHMQHIpNhoA
qpFVXBwAzYyU2dwMlbOAdlZl2R4SKI1qRk7wFuHEtU5Tu66L1PXYFL+vXvzilF0xVxhZgCtGp7/d
vkbN810m4Zmz77pSooEVG9NFFhvvXqsuZdKFSLbqJEmfa3CDu9dBc8TGyPvCDDdlVrEydE859hr4
xshD0+hQdQNUf214zBQavco22bjpb6pM8qnT8bgDhxQYKJBRatjjK6UOn0D1d16j6KMmql6zkXnl
owFHzuKLpjVx4yDT9liH2e73DgLhTgjmd6PkZRiEccTJn69T5NoCingwr/h1LefGsXe3MkA3ILQH
wOV4uvTHxDecxEL0v6EbvB8esup9zmbKfSqTuzQmRR8MuBalJDpl/WLUhfFcvXmdcKgYGl9Vjft/
dO9yLf4ZxBtyG+/+eBwH9bcncmpSu7U00BVn6SDGyYrCVphg6Cd6TFgR2LWX95PFqk5FzuMJidkc
f9SneQ7LY6ugi6b8mCtoWGnscBQL+MZpadtRNi60aFdSRZLUrml0Wfz1hZgrK0smQDVwlyALANW2
+neM2Zs9xFGvUYniRi26KucWvpc8Ffzx5YMnVEepuWo+pLFCkjdi6YYCxmoOiV3EnLZ4wJTf2PiW
KtgS0weOX2sV5tXJAOxVnri53KZVRDZ6uvDK8pAzW8WmbFyBw0OJTlEjtm2q1QX8YcVIkb83mw8s
v88cXuqqdhLRW6+Yxp7dbPFYmMosFUWQxHwZeXaxF0mz2wJdmSMY6McwP2UKICpN6zc464cQoXD/
ub4o65+OOLvvqi+A1fY2VouodS0SrEuxVs4TdCMwzSqu34UWYFoDJO/X266U62VsfGEzY0vqu9n5
tuGKRltKcBEbh1QkVlmr93H8CDDMnT40QQe7KMufiTOSFtywooMrsuqBsWE8wYbzbySZQQsBmTTj
mQ7jxyBTyZDZHqVax16BgJ8HpHwDv1LsTGeJ48wy6FjHrSnYlBn0rbwCcWkbs/NFG+qGny8/U9dt
7ivCh0JWRQAWP3vNGktGjjhYPODRiGM0aYpOHfdJ2KoOWHmE4Bfm1Px6FfwOjbqkZgx16y8qjNwM
k6my3TUpW89QMfu5RMOThE/x2bjqPGYZVo3/oP9me+WwNiTj4eDj4ircxHL/ENEac3ThwzsFm216
4hh4bZVAzNFUkArFDepT1GtXhtk5lIR2Bc5+dG5v4Oyc334rM3qyIWVYE9bsBG6TCOVj27OhJwYB
hg4SVuHi3VO1P5RZqgJtn44aItwsSFyUAVWzTEnNSys0RfK7oOpylwXJJ+7ygygJAsVltV+6nqr7
mFSQQwnVYZiu+soBXp/R0T+qYM4SHUeAXAOOPXEqo3LgSJVCsJj2sWZ4vc6toUY4lAJGyvGaQpYF
174Ra+7kCtw6GXPwEedIJ9OsyPaLMw1JuuiJN/S9hFBF6LTLQJBd8ZoJ4s21O231oLYKLEbvZP4A
oKlRLwqGoOuX1kl86GyV11qKQ0g/Ue+HinOU27pmKa4a5jjq5iCz/dosv1Eb4AyFsxwImCL4D+r/
vateRST6p1o1Zb+Whyvw6Jk7ZALap9g/DJUDIRmdU47oRavGyd4q/MIUGUG/DChZohYainSqjb4V
Oqq7i4HKFXLMFUDZYBDh9rnpyACo3sVVwx8XmcAVDZbiBt9j/DQ4gIAEpFZHNSDC6FUQdcFyIKAO
0d9V0iJq/35eZWsPf3DWrK45DpvBJ/p4kImnJ66ITD/wzoAtNlfZxMkOotn/bnzxQyuNUy77oUiU
9TEhCq/MWMFAED4qSBS7PhUl09pQG2VMMcSluROJGx56JU8oMVdWUBU2u8y0Uk3xWWqGUEr34CuP
4ilcJ7TFIqiYSkw7kxkW10e+XMZwp05EvLs/Ua3pMKkPhou5ma6WlwW3pqBTH+NCxkR0SE/8F268
GlNJxV/6lXXzIKPb/cyb5BpjSpvPg1zKa2FupiGPlRvIozWbAQE7CmqTffMC+erq/a0yUw+30NKJ
nsUguXYdNArome6JbJ/v7eAJz8S6Hkc+bIavqEu6RRoOJE7HIXtYpt7pwsXjTJVEpAWv8uAtt7dQ
BfYoPys1wUmtoXV5k2UHvqRn0geSa1qFHbQIO6FuhR90KBC1gDevRd6F4503f/Aem8wx1ysoOdlT
M4lV9JZJ5vpOwkMF3TFU35X+cJvKW9Vkm1kZz7U6xozVUGZ0npf6NgPvzky9JfralxW6KXKcO1/N
hrDl3bEQCRkdmSAkWCGzkyLNPSSdjKNHi7mJGb2rdj9gQlbvtf0zMIftEC2v3SqDa41bgfZ8o2Ug
B4HD8PQa8qYp+6u9SaHSdX3IQPMm9JXPOCZQKDpwC+1vczbBKjNbiKIPqh7xJHZsYx1RLA8hd8cV
hovL/g+dp6Pr95J6UAnC7qXHZ4f4C4jhsaOGtIpiQ4hEHXgwQE7x/AJ6O7kzN80+xRYh12lMyKyL
0R6Mp5NB0XUYfdQTuwtf2hCpgjcQD3iEdN6W0QP4imlSpm1nnwt7xQFC2rKYvyGbve8Q7pAp+vOo
e7FujaojwvMbelkQNPcBO3jBypsQIzYr+ffkumrePJct+NXnr22CEtiIsOFztWvTdYjM8C0kF9AM
87bBB1SIhnNcqO5BIbCYhertCMJQHD7RnuZ5VG5gJscocfoEohfgaracSrQCozJKxxRNsYBT4uyQ
1+7XVLJmqI8f82mjx6u9LY2GEbpTtfY+iWsDyJVnQRH/N223k0opJiO1SZEKj5PIs7dc9Bc42VO6
rCySAY/xjOArImMAD/V22TLDH+nY240268VsxADASsBeErVux7Isc7Doh+SDzGIU5YFE05ulNcnI
1mATBiw+9Zj4jl+3zM8dpiMuyULEoSdr6jC9hj9/cc47wWOuLFvsNsl3J5zMs8hV3ASZxEReffDN
JsDQe2mK32mIaGNmGeA4YoTOEqtbH1CPSPtWlNEQ91Kvna7zE4/ngRNT1KbMcLG6lCHqpO3Tng+i
Vq9IrJ7JCAMvMNMRvxo/JRmq+eduOfW1cI9KonpjHHZxQuKH9sHtBV+tdFFukN2wrGxpTqKZipmt
DBqkonTHx1fYPHVbfB2OcK0vBVbJEhVu5nWN4OCJ6vt1Pav7EzybC7kGQwZsnzR/Vl/wIyLppAf5
wsYbGAeYy/ml5ftRMA/wQsGbWmOQdNk24W+BTS1+wzOA6OmkDyGGhTn8+ZskPPx5uZW4ieyTArE3
bFR8aK0tlfshIhoP00FrMs6ZmAppxkUxUAdAaDfMl9aojZd00NEDc1+IU1+MMMmtFjaS9+HwO9Mg
HRtwUdEgyy8Css9DUW6TTs5cp8YtdsSY9t/YPSzc82m73J/lZQvxArppSWsxlnjUDKBxXcK/bG+n
OyiZjxy9ajHZSx2KH98UMI4hUmS1ME8R9w5PKtLuwpUcC0xy2+QL+xjDwuKnD+5QcaZo8+ZespcM
BagImeIa0DX6wIuqVti3znfOaccXIeZpKXaEuHsjCq+yWcOoev736OkMBo7ewcMupa6E235HoPDA
5JscgAnE7/o+XEiI8OB55DK3gvb6ibhTMm8bPXPZBvwPG/0Y4osrQuX3MaFSEv94Tmq0sHiDFnUY
ieOGMO0HLQmW8YWgpZ6gQ6jtboIvlkPV3WlhfdhNB9VPinYtDCJxzm7blvTGBGuYbCvyvKV8MAYg
7b1lqbUhKgLEFC5R48FffOkznQhUPj1N0BCtQGjGBw7xjdTO8gj8bv6+EKnSwaRPRoNA/DahBHCg
QukDiLil/unUbn65LVw7xq9QNsRc4vOzSqsxlDZuwG9mtw8EHmiPnMqQYGoVuQc3z6MGNB4i6ZG4
zElVwmQLe7Gtj89HGvg8mnRqA5QRabJi70PGDltUG3lGF45JoplRpJQhdaxojDCVmuxrNs7TlDS2
4fZ7Ls2ZzXWRJjJvl7zSM+86ckkgpnRoL95bV5XwYLPxx1Kzdx470dAJZ7Aw9cuE96eUS6wFwrqz
tte1ESZuSLqsMIe37qu9YNQkDrKzyDRDoctk401dtQnGGo+QkiIR/dmv8mTi1PrDQ9XYxcLIWM70
6l5i8JMYQbdnO8O03a5ExWHl8SmZgZhUS9YNo8ZSPA4r11uK6ZQg8u/quhQJQDyyk5OEgczNG2Xu
bakF088enEW+ahjKt2pxZJQiTbMqX4OjOikSFrM9ROdPNDR6ALDiaYZlHnvsGtWMk4M3NRlroZdE
ZeDiZWkVk0y44ssdQlux8L4LyGe89Um/FLXqFMpIXR059zUgLp+kE5jrUBXKtcOR2+5yh5XC37bU
dBixYNdz0ZmA7etPlAzp6A9yHrNK2BG5d7EctP+Tu67IOhjgQT7QcQPEKkw5B7Gw6Q8z1aaEnv0r
ctju1Pp8D6xTarBXUm+3NGGhWqoZl+jAL6lnierOqoh0e4PvYmfMeiKo7OIVIpZMXsIqwbiFMEpN
Ck9l5L6rlpFj4UeH26Q75r54XWCypuqywm+w5u4P5NFpo6yInRd/AuBh/Vhw5lARzmN4aWcbOi9M
T5rVaUtrWHaf6gLRSMQ+8wPKWaf7wjQXdLw/bk7xrKfyMmOzMfWT4ewtoKuDyXMwRY0NP1sx/aNX
yn5kH5E/twjiOEnOq8/3vZTxFSd+F8swbKhLlrf2DsEdtDIY+zwnACGbEr9MNPDJKEg/QhQbFlyO
e846psVk4OoRjK7SiHhKjbN0lr+q5WKkyzIVzOdRLbkb+EmPBYZ63+oNC95cgTrwsEYPH66gS20g
JKlCc5/u2wL/zt40YUqs9k1jyCUrWuxFWU55idK9CQNczENrirZhqn6IMmGV9U2PyNeZmBgT5RzG
bX4R2YmOe1yj8aK/oMKaed/Eob9yDFdrOrGwyAXa8C1bmvurDTWkqR7o8pL01k4pWpJGzPzaGDeF
lw5dUilOWjgIsBOtRTAdcredLjV7CDg/4W7fGXIx2Uk4soAVXtsylZBvgc+fec/kvzAtODlvukhU
Mc7ndFqb2GSQ9mZxEgUwcesyC4Ahc/x3YbOaw+FO1hsWIOqMc3qN2veEfQ6wbsiwYnvJy1y4K5fP
lj1ab8ZGJGwIcoYqiG5UOR1D+ua/jACfl6eqbyu6b/1hyVSJG2aGaN95pfyk9CZYb665uAsfcPKU
Eh1MbWL61FZAVpcenkaA8o9Y22A8RQ5zoy6kKup5lsTYfSQTE7vPNa37t47npp4H+u2xD/laNnka
jqN8/qIb262r08KfeJJh79YaiNYQNVv2ZQ8Hbnzyx0IRhSMq429It/KVIjM3wx52bN+wf7QqjnMO
3dQeS6YjMuyiknMlUY3D8XjJZlZwAEoUKO9xTIAT2Zkt8zpep4EGWJMtEiFPaK5Gin1IWoON8yUD
2bNNeH1LpQSF2udB6Lhid+nfmOCuCbi8WFcUwrBHiI3mAheWUFFutc6F2kc3zXkUO65E9tTtWhdq
xH695eQAUf+Us22nA825/VI2HsLx0YMUoExJSdIgVZZ5u4EDxcN9S9nfBXgnT0daT5mMQjCGHA9M
e+vN2VMGfC/nmXpn36fgEnwMTsCF7wrLWtoHjN63ncIpuIpUM4NuP6bcNEN/2Mz/ldXlVO/3eKpa
WJeX1nMcNocmqLib+4ZmIakPKaXeZDrcYsIAsGL3rQkhGMcG7Km1A6CC+ReRnny/LW55XjmzXESn
EsZ9/08U+5tOurnNxH6YvL9jrXUmwXLiWyk337dKtbD8dDTmRQekwDmQov29+ZKN2ROFje4czwSw
tJOgtgVJm44/kxB3gY0K49zgart5wUUOld4RtYi5qk4k3KVRqwfyUFBW2H0PIDmipHTmCsLpPEjS
4Lz2wZWTbaikLw0C/wh84dAq0VyUbxbTm7xBWAd6Xd8MDkh5qAGH0/2ZPXK2f0Ar7oaQ7gBBZAYz
QcrxEEogEYqEGPBE5VDBoPqDu6//xQmtj5okHfQXZdTsRV9Zv+1COOXOxKA67q4vzO5ycQ9XghUU
pcfUHUtXeOwAuvrzz2xk4oyMn0eOYRLDY7bmbDKavREyd2lHdPf1jobQ6q0THSgtttsVngmnZ2XI
Buk6Kimtfu3etR37k4LmKqtLtd4THCCHiCsRubag95bt/SZjLCPD2uZlKWHd/MJ/ILMFrPuuq0T2
pViyGcr+7lk7ij6uThlOfRfKMiC3md6WWF0/t2PrKL+otlSoo9JSJvc7zzfnpIdR8wSr8M0HfD/d
WYWmVPsBwwBHg1SaO3cjTvHZ0SKoz7zLaL8rixy+aHMwouHQnVqeJ8pwJ/z2FHzcETQIql1crPxb
+StQpIARdGTYw+ZU3qmH3Ag9SPGz+sqNP109a0DKyw0kvC78W/0UHNewJsiylyI1VeagTeWC1GeH
3d7oiag3A8vuH4KRuvlla4JQh4FeBwiv9UavcPml2PCyMbKFZICXo4eNhHfdNzWoDgQdNedTrCs+
oSrAoe4U0klnyGVxH98xz+00g2w5RhOLaqg4EgyNGpT8rhWGeH5Gbs6Enhz+Oj0w2YDTYobo2YyY
BcpO81lcMBf3uD1hxUtgWfyW/75XK7LFaNputcx9DFKy8c6QyX92ZX+tBwi9HUd9tRdWRRWjBnLd
E2EDUoQKUuWaJiCc388GhxooqqPg0Ebn+8Ihz+v5DDKBcq/U3LcV0+lCNSJmBPjNtAlijrVb56ei
LFv91wjHuoxnhV4vOmJ3Wf3bghcrWSz0aQQvsBjL1TBMNVi+KraPz3R4cva+VSRJ2rTjWyiZVsxs
EAA22ruE7RuK7plM/EmdfEVH7ZxsZDSFvEm76AEdhALTguCjjGpjsyurcHRkKnZXMiyUag7+IQ+n
aSplqZg3xypUZuwTwHTk6xV3nr/WHCq5mNrbZrt/OMOssZQ9qCNjnI8mfW6HFiplliSkNc/49U4X
/uoGSg23YLztCtqznxoxDNRAtvh1eRQvE911mmILrvyS4Pe9RHZq3IlgGTK6IWezKfN+NNIdRCk5
+qVSlZwmcLMRKOuMhDMgFKgd7TXr3UNWdXYyjJvbSIEWx1hoBCOyRs+cfe2EqnB/xXBD7HPu1lq+
Zh1VvnTaoBZKgZaiHdl+7XyYUQKxpzRMzmKgmUOPb0SxEm8z9riSV3fiMSbRG+jajMsfUybNBr65
8vUep8N7WzLdd6ixcrnkeg/fjJVFq/9Z0ntJTXDeh53eBf2u0GIVOsckS67F7vJHMXE/sRORfCut
HmTNgHIKPu172keyd5QjPWi5nWYF2kpR0ySLY436+reiUuHdzxuY67aOSmsgQLcp/N7/TWWrzfN3
oTXOqSoiaWBNXseAXvUW6qKfNrJxZi/IL+HaKGlTGSMWxMhrov03SUdRJmPsFNcuvNTXK40E6dHv
6nkSbijkhRT/ETHPiVG1HvZf23chaN1AfJ5vA30QLi3lCM+HdePSuRSgP+K/8vCEzXpHA8hu35ZV
bCgpJFJ6BZ1qwGzuFWF/URau49VebgNFdSlHSAtY6TF/V7mkjIF3NLO0/eOrzoWhOYRErsUrjvvu
Nx76eyu/bz8fMvHj2GUqRQeawZ7jO0QCiZ2pWAgkcKCBOHPWtu6T9SWHYDZkm1sbXAQtPa0tewdR
RdF+DLR5sI0mJ+91D20Sm3+nH2wsnde28SAXmpIbH3etgQljSVgGnLuNspMRanxlDGjCnf1vrmBP
BkLKVagaWSBA675I3IAaFwFIRcx4T2/e1Ayuaizl1t8s7Z2pOmvinP/JwGXx67Jdqv461hikDc0u
hwzAnFrMfRe6IQaq83XyLDo+03yNC5F1sVP8D9oDzffpJeBIGHNkn/6UX2LBBNzfpB5qzgNKmX/G
PSua4khIAk+yRoY2SDGBS+AXPTNkxGnt52in8QQAldLBGkFBgpI4l4zuBsvWO+HYljaYqFY0EqT/
kXxSJCAtF7lNwoKg8lDUp8r5l8f5gvdKpNWjHWWsPwM4kjbFdTOoTHqXE0p8s6NCnTVL6PffzfV6
CXo6FPwVGo2cJEIkweOuS+uY1HDMP0hhUdOo105iSmQ7UY2Ss++4TeghAAmlDoHdlx3YUuSkM0NN
w27KdoKNELTsn4lhtikncSjvIE/QS24fVZwuNSWwVPjlihsAXdUPcG/1qgu5LryqvBQRlvuuh5MB
DbyWLt2/Vwpxyj1jHR9bMGHdELekqcsSbx/0T/7zgABdQwwM+VhN+7AsYC62dIErJD1tQdmPWxpj
RDqTgsPDpd8brgkttgCtG/6FAr2mkB/q2Z1Yw7z4h2zVe94nSi8gBPb8w32fIFbBKjxJ+P0A1U+4
UtGlbZWoLMSNTlIZprsetvllQJ8UIdmWMoAXWLUQ2nG/3GSyT77CmTLZ2gDxO3a9TEhGeSBQhMwa
fOcSSHoSL+g7a7WT2bo1OFGl+69dZlRkVdBd1YSkA4vub3UXXyDYNzyfWfnSufMm1nOUtNNte5MV
1ioNBQCEko2U9rgcwa0akgZLh3RKH3kLDACNH15MOe7E2dj3JiipBD5yx9sFfklJJjEMybutVql2
uUSK1arjcp3rXghpy+IkAYOQZK/2au9xdYY8n6tCEfRtTRdOOJKgFFA2mAQMx1qpZ00ndh12ENjU
fj2042ZDfTPvi0KuWGClJkggVzCU4ZH23l2OnHssdQtyw7FcwmgNidDr15YAZgDkPYxGuFX4cBrt
CNHwnP9dtrt8XyuNfSd7ffqW+/h1yaS65FavCH+x7O5sZYZfJHmj5QmjxqjeDYdbFxq8PByz6Q2Q
Vtnge6Glg84sZVyqtODwR7l29h9u9Uy1l8rBdtGfVn+j7F+wtKXMnrwP1zCrMyHaFsZQsfHYhl9c
9agQ3rHykaUf7KQNLwYlVD9uhrIG9nAbhbpnhSl81p4vXxEKKvDTYfQxiiVOaSgT6W99thUAmriG
XuCh22cqWGAXsue810Qqj6+rYWcHtGTmHrNAkngJGrVKidIgGZtkgJgvkb1pO+s+pZZaBTTL2iS9
IInboMnDkTeVJjOsEZWQeXTHw2jktrmfRlYeLG5tEv3RgrLVZw5siGlIugj0wjV7jTNWbADfw8RH
meB0nztfDMPVIufjF1iIzQ55ks4cOXjpjBcx22H9Kwiwrpnhrt6aYuDdkNwaIjBqH36NT66o+/wk
rgmOai5nBlqmip+GdXP3RJArQN31GYu+5+sxaDVDMoHqcRXr41BHmyIs2txvP/iQzgfQ1FVlliLs
UQrAoK32DvF+9PsMMqkEGqrhglOkVPtKa3zncT84HtgdYld2wKRC6DRWGjW7Zz13pTyCmQdgqOoK
QBzCYKOWhRMUjqfm0wU4SpxrQTJN4t1GExp3lWLbyu0MEmbCw0zOyCkqqiGAzlVJBzcwlg43AJrd
UQ6qaOy6wM8ERGhy7j2y88lzdfUXKArYjjv8Pi9o1Xvx0n23GjgmHhoJckfp3/YxVJCM64dKha4b
B/UPMYUspAIZt8QpoiuN6xYx2JWbn6Lpu0U2tXveYzKHvka7whIaSTK67e3b/7qcIHIV1ed2FuDU
cp7qKHiUutIzBeXyOQgN+lTLV5nIQNH4wPAEWF9S4/GeM8D68YvD3CtNhSIA9sDxS5C+Z8FJIrxM
IY5TLS8gV21Z99smJAFQXd7fxIJNs3ZLij0YS5eE98hbwL3ertBzjvGvFRB48zSgeSP6Xvohz2Wl
O/vR9Ki6WikgatQHz2YAPjsw0nuTJ2Xr6SHtgfTK55tqQJRwdBdX5JKAmNH2hoF0hqszSuflUdq2
8fN6qf1dwAEkoWU71Gr7av+RsDkENV3gYUHGHAhUeLH0uiGRUP0XFckmTO3UDxaZTKwMkcMND5Uc
zRdb2RDO3N/3/M6+6E2Xh/ukDSNZ53JeB3AmkQhworP8YTDbflsXKkbR13dVrlJG8/tTtcdmMLoV
2nco4N4Vv8rkRE8MyvaasTFxo1XoBopmXiKXAdFFeG1iIufr5F4rFdghKlfhGb6wXswaykZPqUpu
3kE8o57KYX0UYJ5zV7BM2AnKLg1nzlaCIPR01m98AjrHItm8PfDHZy0QfBxuBXr6/mGPBuCdRNSR
OvbqD5wCjcFD7CCDHowUpsjaAc/d9kCuE0yX21qFwqXLnml/AMItfZUuAr3DyK+kqzIpafjzoHtR
h/EDcwbokjPav9SNJN2eqfoM1SiVV+5OXH5ecVRvFQIKwtXA7PNrfyTuhkXxYkvzT1xDUFS2WNfa
FrR29xjS1H+cCE2usDfvceQaExZwAjfpmrZRy5EII/OvgBCAgkfJF4qgJ4p0/5+Ezv0EkWKBC/Et
ZYhGiYJTpXWrw1w/qc+JUREBNrx9WI7Gw+fOjlrsmtQDhBA/z95p1AqpYE8Q6P9GEgpfUEbkxkso
9mpvaFP2GhCLuL6j+0Vw7sCnb0H4Suk3E+PXjtHwiWTGgCLUO1DQw1pb+fWB4cu8jTX4iajaZR/k
WmWg0/hXULjGXxUHyzVCKLQ4B77Mu81Year8VwXEutDs+DTRIJVOPFyQt5yzbx1P5rD+Q5zyoDmr
CsJUef4m/bqWdYy4hVU4ZVgN7sW/fhindRG3fb2OiaD49O7Bx3jyTy22w8gv7G3Kpl+z9jYdwlS5
ftj2gU3gvWkOaQTU+heHhn39g7Blsjh50PNZpp4XWO276XvNANxCDYPSP4hlzUiVKTwlrWq0GlCd
X7lwN66gHM0CJF46pWy0N4zEgXSC0rRitZkiYPTV8zM3YBnFV6/8GD/GB1GXMQBTGjCWyZsZTQBd
/XZUsRlwtPorc7fFXZ/eIJ9oaJw5CE0X0Vp/CZUHQU6rlwX5BWDUGKkwGlzSKoqPL11stFbm7ERl
vMu4wTYlkvXHimyk85/M3hZ45SlM4Uv+Yu6fWG7zVcwZ4bgBr+Ynf0380mbPUUUt54tqy06JTLZe
tyBy+zYx8pTRHJD+ExyBnLgzs/IxPA6mKo5Mtjq6rpmxLMs1fGNLI/mAe9yKJi96pgwZWbvH/KAT
wKdraEDQpk5VJnde0C7nmz4cMqP3NGdMyh71SAH4bd0l/HkqqqW1hoKB9oVXDk2hFuCINFVHFLiR
ZretNZ8UjvFkQ11sE9/c61HxoRYdlLxwZ0EfF1ZtKorfWDjj4iB6aOIAQseS7aNVMHuzMpYFOGLx
iknc4Fd/YjuzVgviSyVUUEulcBqkpwidFNVqx1EY4nwWHh24Su37twhWRRO9WbT4IwqfNXNuS6cp
ZaoZ1KeDmM/MYXpghldxMCsqkHdXCc/JR5GSqf0IpPVp3cRLyCpQDQ4p3TJzWV0NyaQK+5sB8h3v
32ryyBPVglWbADyXGzFYiM5eQZiAXuCX6RdJrZJpzQMMD367oVsYx8Q7Ua2MHgR2aqheqZx0O7RT
bjgEpZkjCOA0UyrDRG7fkAB89t4ACSz2brN22Kp0GMtjKoj869AU4WRB1BbL4oA55QCEAssZ2vPK
Z/N/GSHWvdJh5xk53HLWE8adyOHKMCyvIN8v4dFJnlS8j1XqFd3CFYSJFkPjZMENqPAiYpKCxZKS
SzksdXn6TgtWTY+moSkHyjkfhUXJ5dpaeKZyJXTJPn8QgGFJjJiEpTt2+DmOXaftXe43AyEZaA2e
ER4OnodElLgtOdiXaxo0dfIO7SyukokWHCFTNtrNuj2kUYrlXbwo/cEwtV1nIXFQVBaL3j1jmzBe
SJ8lhOUc3HANfnIgCVO7NYRStAacCI6SGni1Kpm98YMffnevXeF0Vv9bBfS/CFKO0Ivy22geRf2Z
PQC2NpUww1jy+VjjUCYql8Z9Y0xY14ooAJD9XE/zqTtDv+tPq7Ch0+WYHwgKr0dioqb/0JL8D535
FruSIoRpVspzk9Du09JZOyVV3ZqZcU+8vN5Z6/qwJGUGUtPZ+eWFZA0/tEiKoDc50AfQpweFxMgU
YcWdo9+XDOu2l0FhsObETWWsLaWKvdZUSpIdhG0A+kHLJkDuIB9oJliN9jIyZQbiQd9DgDnQT8GV
aHD/JpZMI4lZse5Vk/4H6FVomzmm31Z8RSTRkqIBponsMJNpQhTXqQDB2i6+PcYlmf8eHbbb5PXl
JTmYd52GI3AAqAPXc9dK7ehlVrJmMbsPNPWxnZa0AMR8qy8nXcIqYZDOxeZF6vwmpm8oKuRATjXF
W5DT4rwzgQkuw/invIW2MoXd4XPvCQQfNJ64RSnH3TrGWA/CNqth24c6+BuhNby7YnAeIRP6oxks
19dWQyx6sqw44dUpIQlQdCrDKKCrE4la7a8jklTPL7Tf8Jsjef1GbP8vyg==
`protect end_protected
