��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����N~@#�k�0!����+��=L���0�ԴZ�2�Mc���ZO�����=�����վ�	"cqw��a��TS[��{=:�����K��-�մ�(��k��N�-� 偙O��QZ��~rL'�x[�i,mׇp���O�I43��4d�,�H�����SN��d���3���r��m���̨T�I;uj2Y� Er�*p�Q$Gm���p�V�`�2^���,hz�<p��l�Bxt�5��s��\yq���#�@W���f:m��T�	,*�񞭋����_��㧋l�	�\�:��uGd��PǷ��N�I��_����Tuv� ���us�(H�~�{2H�:Zor�Q	#%�3ˠ!��iS��95�,?�.���/�F�i{#���Tp5����Ҥ0{%���2vpn���X�����@l����3dc�ק�3	�Ed&3�ZN O���z��s�yxӡt��v*}ԫy nj#��lc��m戭k[��5)�A#�����8�!�]�Z�s�M���t��w�!��'ÒE�rv��Ϝ�c@<U��\tq+��&|�&X1)C�����r�A~��B�&�����s�:n{p��͠R�X⺂L^��R����c���f��J^?��ܣR�O 1�rV���:��T�4���AD����˩�F�w��)Dm�O�b,�a���1$��c��7t[i2>�ޔ0,S���󧇳Ϟ�ᒨ�-��}�!6��Jyv�醊�^_�(�H�(y^����o#����X��3-�k\8�M�T�"`R�DF6ȕ� �,5�;Ҭ C�k���1\������k�t־9�}���� ���QHF��"��t�9 ?��{E_�7��!����](�S��0�q��w�9��=�i]�1�GʦȪc�W�XC�|�$��}q�6�H��Sy����=W��T�lêL7�6��">]�q��U&�,�x���v�5n>K��z�b�ȡ6�a駓�n�|��W͊�2 �5��Nf��5-@!3??)�?&􅣨ZT�xz����ari'�ǫ��;����ȃAw�1�#��(6(��^r$ܪ�O���3��4�)��G_�8�I�g�(�x
N��C���Q<:�]�BvOK�ŵ���G�_�Y��
W��fzu����z&I��۳AfO�B���bhZ "�ɸ@ .�Q�H��P,�R+n?�I~2�xN�ՏL�I\QԵ<Z����`�擬/���;����ȗ��Wx�.����>���
�+zjl�L0�%Y�D���Ԁ3�xC�^�3l���©e���DqG;�Z��;��������`f���rckK��ͼr�+ �?�A�4o�뎉����&[�Q0
gը�`��C�Yɠ�
ٍ"�n:r�g�}13^������I�*�K��>�Zڰ��ב`*��'b1h�@� ��h�%��(����͎>��5#�\v!K?3@��K;P����qh}3SZ�P�ĵu������
	z�gّ�,t?�c*S��R'൤�]W��KC$��4���14(�|��?dY���o��f���=�5�:�u���ɪbU /��J0s>���?q,�l3���S)-���h�}"ZV�f��-����yWMy�#���ȵ����

�#-����E�^d@�[�S9N��ڎ{�y!����s�@�/���õ��pa�:Ӓ�2\7(D��S��~f܌3�|%�]��ֽ���^��j�����)Y��U45�r���
����ƅ��;]:�\?�� �����2��>#:�9*�_�Wc���� ygqU��o�m{��>ڙ�;~��u�n�ɞ�Q��r��e�'�'����M��{i� ����{R�c�g+rN�]-���L��" ;�w��Đ$?PC�q⿙ӿ��;��f�Li%O��<�$@kK45��2��_ta�O�Th��q�*;���j^���*O�2���|��|�=�{>Cf�8MB"����&�yg z�໫���Պh�c$��w���`�C�מL�����S/����F�W��;���Pm�:Jem��b𧻓F��:��B�MJED��s���Y#�j=�b����	kb�4)��%�G��NW�(z}���g�M]����1��fvj�q\��?����j��>�ǽ3?�l=!�w��X�����=x�)SXz�HQ��Yeu~�O��Fxjެ������H¾�48πwZ���(�-�����������Y�ʦ����4;ne�D������@���\-}�g�q�x*p�v3�a\�;\�Ü�?qw�ہ��P�q>������v8psњd�s��Q
�FP1�)8;��Gh��_���cWC	�z!�\s��l��5�ּ]��_��F��qA�78v�J�A�by28��1��	ʐz���uj9�d��{��P����]�!���pjCMu8t �͵��*�����P..qD��]��E����R��ԍ%�쮣�E�q2���]�r�I(�&��q+���8_�k��U6��@��?C��cj�_��k�����oG�o)o�J��F1밒f�T-XP�m4fd�Ȅi��Hj\���Qz���V>z�b.�	����L4���^L�%A��B��eK̯÷�0����@Z	����mr�)��t.R���dQ�_�7�LiG>]�?��ZY`Y���Tθs����3W+@��71V�Q@�[�[�L��9�/c��<��mR�eQ�R�=|v����\:W�quD6\u0zj�W�x�g��{����t��j�St;�4�j�K� !�O� ��H~*zĝ���H c�ۭф�3�'{t��ɢp�NB6��N$��m� �P�ى708+�H۫�$
��Ip��<�͵�=ap�Y3Wq��Na1���A��`�'��H��>��[h�˄�����3�zZ�=���?^I� �Ú��<��޿�-s�Ū�n��t�̚!b��DL�i<�����e0ʊO����\����}�=N�Nk�}��\���<�Q'�jK���`�	���W�r/�Ҡ+���ӳ.���[�>!�O���ӬJ�zP_9��PëZ.̝�
��?��?W�7�~�%�e�6#�-��Ӣ�s3��^Y�|������0��m��Yx��(_
�[Y1�>����l��;�G0;%�ݠ\U��;���c�d��R2�4�i
��L1�����bCOk�^�.(���z*�Կ���FN�'.N3a3o��MՋ����ģ<ڨ��Mr �o���Qjw \���j��,Ӑ�,A'F�a��A�<��r����������2����
��?rzpռ����e�MA�k@^Ux�e�/K�jHaA���,%GHN��hس|����^9l	y�u0$�r�}��q +��(e�] Đ�~�M�}��Y Ȳ��u��,N
��fw�Iқ�������_�h�*gnJ�7oG�f
^3�F�,�@��Б����"�*�{��ֆAmٺHAЋXȢ*��`6�Qz#��g*�t�����Ӏi��mB9mphî�I�ͿG�	�
/�bY�۸>��ȚVg�ݯ����M���,��fj_U@�H����\�s^ �5��bK�m"O��#2g�,��Bw{Vg�%-,Fv�"K��P�a��Q�Δ ���6?�jM�K�UbM#�����>�yq���N'
^�����-�,6C�{���!��< �AUW ,��ݹ~yI1Wl)S� ��W}7���D�
�n����_�n׷�H�mPė