-- (C) 2001-2016 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
koufcR29hJVdL33CDWaySsYMLKvWsF3jcTOiF284SK2TWsvUoJbDdPqg0DhvJVfXMhduYAwBCsGM
dPoqw2IIY/9y+DOmHGWSG5kpRp0E3r8DpOndQhB7sXQbdtIR2Wydrt3pHdDrqGyNy1zZXkdoBfQ3
y5lD2KqqwWQGOFAALt5TGCfDMhbbshlt7adKVivpQZ9ntpA+NSKsl3M6pD/acT2wW+uIXiAWZqwt
iWuJAJW4R0bob5fB6X+iuEIUAEuUCIiDQ+NQGhu976yxhToN8t9wRwZvuhQOc7LvHnZiRXoTRX6q
GCWUbNX5RCrxKRhffs3pO8oYXpPVUvpJM0Wphg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 4160)
`protect data_block
Z1l4AkvJieXrlTEWWLMNN3MtYg+3dJqjU9XToFN3oQ/oNPURHBhSv0TmOTBQYDHK37tp2VixZGpd
GQVDm2b/jGIbGrnFzskWhSWP+9GFDklW1nGrwhqlq24/U2VnAye7xDUMiMgaNXncKJFfR0GAro+V
2tB+v92nki+JkIY7Jb9VcsJDcGWHp5GCxabbpydzxyfK2ud04PbFYCouoaqrrKRbmZ2ECxDftMBS
SMSNNKXR78pC77spx5IoV3TJDDjc/greyE/lfE9WPX/e3rpckb4GjehtNkwf2Cua3na7mm4FFXWi
qRI5xcj8QkEf7zZ8MkubP7nIU0EFCkuVnr3hQhKeoT8IXZKUlFPgd14/N7WWUj63lKpMQwMIQj+c
7S4BVhBWT3jQOpw1LbJ9DdCrZePI4HpQv8cVECksfU8/mRx2DaCVpKUaAu6rbMD+Jze7oTO/Zbqs
9ZdCh0S1eUlx3JIGaf6Hbuq+nVGIEaSh/Ai5mZzU82dNFMGkdnM5qnU5vuv/UUMyF+hj+05riDZF
2ax5spGkzh8PdSk58deCxEIsc1L28y5942HdaXY6+mcDb8rui/wgqLrv9+YyJB/YLDHev6BYFBMK
CwKF5CNj7srOxaCvvwNCpwUGadU/ESnIjkMq8aMy0h2vy0X4UAz8Q3nSFjB2hvp/PnEbpYoMcIaO
Yr3ezqqjnv8b0522AezdRSHwe5fLeygc5nY9Ldyuzop4pDNVAKZXTYzSUeZgHm815aTh1pCYz25l
ZxqyAFcuYs1ZiOSTPayK1UUgsnz4jImECARcH0mGXA56gKeDDHQWc2/d9uadKId7sbTMxDp3WtYU
p8+1IqPzANqYBwHCiVxyt2XcBKhHByjIZbFrb2WkrnVsp0Pv7m3jT46QJaxSIUHQcmhZzwIXJfxq
2rUJWvoS1XuR6IKFdjjyfCWoW2UAnFQ6psF/jkhAfBBKapclmbQmBUCDcF0kmGBkOqBBctchJuAi
4hGpLxp4yJ2cdNc1T2TDmbmfzWybHsEkBWQ7xTPje+CIjRKL9qsfQ6ZLiCJSeQJDLCxHIZYPKgTV
LKdEw45aUpyOvcFXgYouAx0IOrPIVvAKAqNGrQGcAiPLqTk/I46F9AXmMkXk1GjuMlIjb8JiEszE
zEtwoXo94lOwwqojLhjkxI2x9l4/zEXrVAg6Hj/fnkhXycwwfAJW7YmCxAPlWrgJb93dLBMreUX5
PHIYlaS4RxBtieIkn1zWbr9v1KRj0rBFI5Wrh+syAu8fz5bH/AoVS5z2WDjuyKD0UG/HAQc9bu8c
LIJzfXJ55OYnu2FL8cNaaBB727Rgm9rsyyJs9IZRxr8DKgF54S9pFgbge7zpPDqe+vfaz/biaxP0
eLtH6DlVFRvHnt9pzXCYHfsSiklOgMPI6g7zaEk2XkKrZ1w1cJCtQ5LT2MOi2ITFriAjOKxJMEVS
9XPeYdTteUDrIM5I6+cXq4kSc9Zh9r9jGeU8Sw6oyAq6VnM3kvgkdNAcRcUuoXJ7T5BgTJ6qD2pC
ypVICIxwG0bDC4taPc2yIRUr70Ekfm4OSahxrrz8McciFJlAosylLJPmujXkJ/7AhvU8eWN1pCMR
i3mfdUZOOP3J/4td6iO05Hy7/H/qoYunF+yfK23h6oniZ3pbE2kOzNu71SHswYZO6XpAWuYVS9AE
rq5HyXWbBTMoaOTW9Y6F2uVaLgpmag3Z7VczCMYBIRUfu2HRAO/TF2oSUGSkDyjEsz5LBmce2ozX
r8e5hBRfmERlQ+BatZiyRIssZMkJ6kcfMCzvykfTp7o8dIh5T5hTdlPbk1dDWOehSQbUYdlycRdj
/1FTfA/+YxeHnRjqs/MpmL5yrdeItU6HEYCwgHX8qzn0KSQfSVztnFIix9sw+bKAlRCG1HiyDbxD
2V2ONzBYsXfbqrNUrMdyA69FAa2jLfWK/qDas6/zIFrKkupNHFcmRhid3FvKAUh0JfvbMKlFNUNc
q1rpeT5XfLEhmZzskMyIPZtNb8Vrh70Xr4OVAMcctKAiVIIwGMVXCUg54UrnzCJALRUAFLbC27la
cGhq7p20Y0UvYhk338BGXPYrGDT+KcPSx+KAaV4G1geax0OsfwQZpZtELRGpEpagw4xZCKKHzD2L
y8RVtV/eLebvqPCqHrTUZHWkbLBQeVo+Y5ZXa0SgTcNCLnDBSYQegErm1G8w8zm/Gjzz6OyUil9/
CopHKPrIe6xukTjLvHzUxUX7LqmBI2/K1TbBKCF6yH+2OhNjfJF/N59A5O012yUTjExtqlWi6JIU
De+wKmbQ2pXeDvtHgh/WVy4JoIn7b5V5GaO2djOLJIBknNWUuRGWEfoYUQ8cTh+Mi8HJmLrBdasO
ZDGVEq4RgpWVugQ1XMPPOM+Jmb0VLCjHaJwu3uDGkca9rxHPyVdZu7bcY2EhckcyymLeljszWzfL
pmjrJT2MeHg2SZTyy2dJqDXGqjG7jhBx3GmNcarVD+m7TtV7xGXTeMd8syFCntdhOuxF1W6RufNr
r3WhMtutDZbeQQUJfrfOqSLKLaZt2owVO9yg2fgkq31ESGVqfqKNnl+0t5o+Pg8Fbw4COKPFZ/H2
ZhjzHo30rEtj1FOBrVWOPHOLlCYgvoWJngjR2MuN+KJ7cdRyKC2vnOLKL3Dsvp9h/JXQS4NJmPCE
lovt7KQgb6bIBdPX/rrPTF9apP7kydUHzc6dpRs3BOwE+cfYQn3ow16V0RWGZXYuPUK3dvo5jedn
qtW5W6ubE7bSFaJcBMOfdQA/BsWzmF6rUBjkL/7jrkP8wRhj2s1rh7qL/ycUkFgNrUgT2KBVir0A
JqS1M/9ZQUnYkfdmv3RcaL2461/6bcFde5VJbx+fKpQm7Q3gRoB+fIshIHd3YpDhOtYIxJAlODBk
oAW6ZRG3wS6mxbEeIyygaGR6ojqtuzaZ9bz3rwlMUFx9x2znsFmMzNRibbtz3/vqtH40puRVnbmq
9kNxdUwq2Z6LZy3eVZ+10bkcoghttvdECweeoP2ZxNOgZVEQKf1IidqyGjfb6y2FvsaWFK0NVSKW
2zqozZ3cTPNuEoH55WC1cE5TcCBc7Ghusua0nyhvJhv9+J9NZdCDNVigPjgDyLsgqlf/09rp++qK
xy85ByfE90ohwIA0ohB6q1y0vvGZIfVgG9ATnH0hUtp13xlrNSrK9xyw7Y0IQES5G4Fn/LvHRzCn
t8WdloMPCrv9pzhzDQpLQxqZoh/7X4+RnEoUASmKWGDzFN5hDbPhDNevZ3j8oelx75YNpQZOBq7p
HqZcHB2oAw+m3RoIz5/kFF0ow44m1QKnuCj2MF9I2wuI8sCzmyxKp2Hd4m8fvJVNxURXTXLnWY7J
JJ9FB0O9OvkkRR+koYvYrDPIVytRz3Y6wDz5TacjkAcq3we0WDuFFIMZpw6/sHsDprEJiDRzY6L8
3RxsArUyhOlT+q2xuVJuvUNMFe6CdjCO4t6wMq8ujdjsmB7TPqRswgt5DXjWC75AOcc4ZWMiLG87
hPhgcg9EjV1kCNSgUSPIjF1AZpdnuRUN31GzA8/qWvnNi0ynvUeIwZVxzzJgzxyQbIurqdtrO1Sw
XRmSV+PDQPeQpTAewQGU0sFkpGPgP0nKdDgYqJF60yZ9YGRbOSdVcICYdzbyqR/OH1lC85om+dOf
8bh+biYrS5Gh589YppDfRVzLThA+ZaB9zeETvlvP2OoEdS6czAdT09ZCy5l4Hcm+RIFoM9zgSLDE
9t4QZFDeLV0hD12UsYzDccR8pU2Dmm7mOHUWSFJfl3LhBnYx8Vt1VM1Vmv8vHApYDBJX+taKh1Eq
o4FO2bHwq1tGwpjEvKGV04EoeVLExc6GTO0Yyaf/cjAjQA9DgchfaP6azNRlEpnhZUXnJtoui6G+
5d0LWfOxsOfbb2qBwxDC4iMHq2PIp0m7D5rUPbS8ZYj2pDgY1XgGa0oE2PjnBeqgKrW88y9vK5Ot
Kz9op+E6fe/xiwIHcINaIeg/dyzvGWAcq2/T3M+ar/fijcqF0wB3KEG8tCl3gsRdYvXgyWOXxOL8
7Er8VJYjsmUos90kXagvCAg6xzkL1P2BZEeUnMvdr9LQodrYUMsbQ/My48T4Gl++J9SSZJkw0AnY
zTvBMJ4CkuEc1mpfn+p0VSHr3yYtK/L08PEvhAeHM5Cc9UJVcClxJ/08I+m7OsG0sv6tYM3iPuzu
UztutwbbsUgXQ84nI7Apu8GnG+9D/nshEcT73iqodn7e1HAd2wVWhG7vBwxFjecQdRNXeELzVhOC
xVR5Hfv/Abe+4+eMqz9Fpz8W2xkvO3SDDctaRUR7G+wg6M+Bqyy7xQGeHfMIrdeqFo9igBPMlrDK
RszlK8Cb+NOUTz7rUGtrmIZGU8bu+IdeRtol1f7RSyWWoCNio9E8qSia+CZ27DthDtJwrD652IhL
2r2G+vMFhIUkR5IM4vxUvAZRkTiWsAskBppqNk1Zfo09mpnAzZXNwxmxa3bIDCrL9GiUFGBf9/Ol
Lcg802csKQ3XbEXH2IsMZNQTsy+wWDWEYvltNPiQqyWo2MVsyGrPZsUKKvccjdqijh1yuWJWLrTL
hIS0hjlSy2r76DQ4tcAWXoh5vo2FmtbZgbfLUX9RraE6U0LHANAjeoMCbkMjUeqwwVngVrAcop4o
0kG3Iu5wahx14E1wot8DNSKaKebeLPX7sBkRYT10Xz5ufQBaLzGn3wEYklkkSxxiA/EjZFj5eKM8
Uinm8d0tT4Jf85wP6qrWRTPZIFjBnfGW3xpf2Zd0E7yQY55ZIxGD4N8oa6N8C0PAY3JM2b8S+SjM
AE4TFY0g9fMmutuwU9RoUMEEajSLbPXULzC1yFwLiUolKQgUkUTOMM2k/pTiF4HFLWXJK9VxGUo7
JaDRbVU3SooyqF5A55DL+GtNHupPeI1i86bGr+S+EEFKT7/csCyqjbXLCcW+bmgVu/I+SCp8Nn8h
tJ0eKJea3YAKZgl6LwOSMsaZgF7YgAe87bnGQdvxfSJaLMHO/GcfcaC6gCDKSHy3aEiMIiMM28Th
aYJwp1ie+hC82Zfh63QPuI6hZVdL5knOF8D+VA4uzXLs1KpTWPpYk+55hUbp8ezwAPbji8mJfE8a
pgYuSBtFDkoj9OSbDfszsPm6Sl/rvVWCl8cfdCR9EAaA8+wByMmD9CULe5B09BhTEFXLskYXVr3S
BjgZzs2Em+sLM0M1bGr25oQMRoe/vVoYtg2zFDhTFetgsKHcgmZnn8DzSfkPbRNJgkh4dd9NXFtQ
abxMj69bbCnrXWOu8yux9Gqm32rhc7oHTga/7VLeHcKC9VICBortYkIymGgplpbDBH6rdeodlMAF
XJNiSrGiLKzF8GYi2kXr1boTyrTIDLgf8TDbeHs/aywIfbXfigfVQ7yIVxBmYMMG+30r16HP99cU
/GaLQ6BSSeq1XQ5tXUOBNKsyVubRxAiANW2Cj1fmAMrrOOyR3RC1jBcWKoCcmCeBz7rhl9MCgAFq
E7mFd4aQkujGRfSVUmoBkSv4BNCWNW0LdyTzwrGUO8bK5X6QYWApO9I57tHsn5TosMQv0y0T7LM=
`protect end_protected
