// (C) 2001-2016 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
IXwxsMmZfqcHc4NYJvr3r68gKpH5T2jnpcb3m1J7tg3XCZwvTmCm6h0hAy0DBqmg7vHWN67b3F9Q
LdBt68Pac8SJ3ES3mSFXvgVBxpHKfpOSF3CCSb+y+vqMfoQjbYWpn3WgRU9XNGAbksDsPbEuY+Q1
vmwILCEwDJnWU/+kQRJwSV5JRvxdzZOn3dDfDJAobLZNW1Xx+63pKISSTaRdkIh4WvrDcp5nNTsh
5Gj/Q3hkj/gxBo/39jHZ24rcLfk7Z0dnlf/AC+6TWqHzzTNZx1VsenWj2lH3+sfWiS+9j8Zrj2sK
izIQ990Eu5weEwv++UXX8FHOYDau3HToXDdEXA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 15152)
AEK1XnW3ACyhqF9BdtycHL6dw43vvGlIvUY1nEpLMkpDJWMHNs59SeY8GJjKqwvhpvsn0yUkdvzY
Vf2jMY74s/IShFhvXql5hKKhPu6ZhoCaI9hXnyQWne8rKOP4izTVnlUUpfCisfQJEz76zo/2Tea3
ZK6MH9FhmkuDI/2snITl6wU5Tig5Ow0+nLyMOkIMSFSgMh73hL+U8YycM2QpEWzHrTNv8E6eiNIw
q2tYlijN40ST4Jq28Yu6z8b3xQOSTwRxbraCgMZ94mWcDrBfJ5+U/W6oDzgLzVvY6LxtiQ0O1RGL
Tb/muRmN30DSSDxJdzSWCAFK03ZRgV7Fzj0DWOmTwVtPqnf68ktc6UhULwRlImLcdt8ZKnwjUmiL
2wS6GsxVRVd+hz+m1b/YqIejF09JszR6QqH431AWAgkkwK+cspn1ysCK5uZGfgWAUVBJKfWb5YVy
l1DooN1162OdMpaSD6hWwKfnvGp1y3qGOywK5qiHj4Pzh4aGrLTgV12RtWvZrY3z2PyMtB0FYb9D
8rti0c0SJpLG6Jm9btYibt0VFzCQVfmNXE5N9NjYSPORdeAFOvjeCzxY4CHTz15cJYbO0XUotxpS
YuufpRmc92V0STn0rjGxy6Z9Hes2P2JaZtvQeyT9ULDpLSL1Zfmp7D7yepdryVR+pJPggegE3xXn
a7gyDqWI1nwzGFh+8DOI7oXR/Wa7+F1h3hkMFij8XXyP9pSoJp1w9xmmFbKNE7V5ib/6zVSifI/c
f9yhSWCT984Df8LFZtBBi0hJa4UVL/RCfCwcrJWAmUYOtK7XEyKDmR2Cppd4rWzwef/uznP9YiHj
hCiPDbJRST8EEOB3fCCJ4J+GEiuZAPcEbgNRfXkzyhTHAMWlHsNpWpU7c8NHVLzlzh3H910j47OU
VueZpV2ezMEPsxTMwQ8MbI/ger9hZ/jYLt2QG+q2IO2xUjIPaUPh2WZ4lVYVbvPLPSCSW7f5LTh5
HixBv32KL/Yqx8gaiO2wR1JYcjMSGl4v7gqqKWjxyh0t8dA3NZhDxjesMhCjy33H7XUgI7m+XuBe
EeUVfno54DGH0Y5y8Oh9yvjexMQ5ir7ArDGc7eQVxuyyxACC8hlX8n0dK8E/gJar7oprX0+kZsQD
cQamjBdFT6W0nJs4T6+qmKDNWFDzrftABJH+JlTidyinLU1Kx80D9ao38/37NrYBJ8a0QCSMbygd
smQIDft+E9Es1bO7F2OTXQVoUo660XkAp6NTRcMgjTITPOxpmNDQk0vSjBBK8CEX3rIoUb3lbqbJ
aUY5qpvvZXR2UkrxX61yHuTdIa9eUpiHuDBTEBU8obdZegKaG86HHmtLJAtEEKfHIwLUjh7SR+ct
FOpxm4UA5oE/6Ir7tXo0bbDm/Ow7jLcnggyEE5Zv54vedgn68Uifans1fvdM3K4GVhviYqN+c+EP
q7kiZ0eSMKKIXO776f4F/N0geGm4yzYbCqNl/YlzYcbPf45Iu1oCDB+gCGbk1xLW6aOJVY5nD3i9
q0vdDxzFbDKKoRS/Bpoq0VLzsSb5GVJ8/an2U7YuDlg1tt7VeDmkzCUlCZEUBQ3g1kJFxNJt2hUn
JN5mCAt739QLjBlO7RD9qiktoVHpnX1vN+UTqGKWN++QFh41f8VlobFC3UBaeXOMKSpKbdib0Bcm
HSZSZYKZOcdpOI6PxNWChW74v7MYg90TXTfns5uETWD5MjQ2zpQ3arRRoH7EfgeABBLzpJCHXTdv
MsQlleYrcf8UM9XsJkscWKiYBEUKAEb1pS20/Onzw89KhpOEnAM3tMBtj0/6LbOeYN1gV6uRpGKa
uDfCTZhC2Amyvb7OMjoCh7dHbe11SFiKGi5bIBYwhNL+53dFw6N2tnBfyfo/HdDQscNWhpuhGviJ
2LFXH512B9I1aNdj6o+3oX6IQY8KYt2MBiHX3s6T/HHjKIIUnh+T6a4MGIV+66hA5m98/gSKHPCV
X+kg09BuB+lY5eackccBGOGI2AbzPglalFCqQMOpTy3QW3fdbMZZ1IkRJ+99uaUZOSwI+uYL9rJD
bf4kS2sqOImHVNriw0wZJQeFtheCS2gOrzep9ljdvoVy6o7QU87GCwdObS9NcdjuqvYwZRpwy6if
vOfTqtnl2syX55I5b6hEx5PEO9m5yoYhSwarTrze7GK7al6bLHO2EH8PCXiccK5NdObNZm3dINgo
M5Ls1qXlG8VClv083AwQ8eCoV0Nd4dL/1RYAe97FL+mawypUe0H61RZLuuxH+NvvEEnOyeLILnzv
tZiid2Pd+WbULtUNK5mF2y9h7PeyutfzihGcXVEgWLF2NzadyMQdcq+rPTDigwDaxz6hvZRCa09L
dQNoxORtmMBibG6tnF2NnZ9HNwhR0CsHOtutIGs7TxEexOrpdmIISWvJppSPnZR9yru5DfWjXT+8
Y6IP2PaopdCCDA15ns3Eq8FKjZ09iwLYNP9fX4NsMn+HLPyzzztg1chCc96+XfjKByvb1nja78/k
t1123cVANZuefjxPo7GAtwROJhqhVLYmEfvhk+8r+vdQYf1R0uHdY9z/1xVSL5vS4pDUA6UlCi/n
ZSioBGsmrTWI5HSqik5yCtrfHYreq0vgeKaLU+y/cKl3PSedg6FF/CWRafm3bb9Bod38vkBWM6VD
eFTBUanoRnjKRRU7MH3iNVaJ4t2SbTSklmTIvPhfkgVCU0MPempLPGRnt+cQyyq3DDf+pLnfVnpB
ewA9ZJFIu4crypN5UQ8sa/FPcD6Ohgl3mlItUG65/JrfwcWsoGStJMWScaUuIioQFUVG7LXo4DAc
KQ9ngFb+mLbrR/lhZNPIHN58s+ysl4RU1W/v7VbsZh/RzJU3PmEUiUqduNgoAuaqOhZOr7HGhFja
f4hVurMcRWQTD+TNmQxyhWP8I3ARhoxfVaDecRmK0Pzp81VBI/vGf4R+j9TmAaLjUhMiSigp3yBV
w+gVTQ0O//nGrN7Mf7K4wPMkbOJ9r6sFN0jibTs56Rcwufb2946eSVFCYS6CcfK0Fpsxk+nBl8fD
x/rn59S2juw5pKv0EOzioVbve9++zlv/ObOjj+KSDx7Yi2PmDBzVIEmZH9W8Hb2vszcGjK6gEpnC
RoptwkJZnXsB8wiokBPvaSwqUYg0oE3nFF1RYet4rnqTaIAmV+4mbtU/oxVkFVGMsMiWrdKMMqrr
FDt/98BcJP4MmTF2hfZKLuSTn/pwJizxkyPoD8N7TZZHYOLas1YzCi3rZM2ZlGwzdSiY77vgaUiB
y3jq2Vg65EVLnhz5gQv7E3e1hCWtQHbTObPdL2h0po78yxSTekkLxXqj6QkgXk7Ndt1PdI9KU0iH
pAvIt4qP4kvDNS/ATiBOJmiIzPgK5TNAduaOQMwjfbjMIjImft553NPTu4dSavxvUpzXbNj/52F1
ZidXxs5NtTg1cG4V8/c1Dl4x8A3ypgVIrqi/QXM4ixW1oWp4vEHTz+d32PsgRCmtQXE7WwrU9uQC
CSqeNb13iu27kbBd7WpU316vADhzLkjqpcgx+1yu4ty0j6A7MhC3yrD+4vWwG4uaz/j7GIVmB6cM
8vWDpOP5F16C2Cd1lCtDyxZpyJpXBQlzJwwrMY9u/Dx2hazMaDWx7RLxR/98TQJsDp9VTgOeUZ57
JRlsb0BlDHX25dLab50SbCuMCINyNqnkS4Xuk1oRMHccXfI7I4EBtT3cYPRLLW/BuDwHiuYJaJ1r
OsBLTNWQXKa1s5cOvMgJ8LgkkvFyQH4AX4ybdliAZd1ONUfQpYFwj7B2LpLRd5PeVPRgVPZwbA3G
rZn8MYg4gt5qyk65zMDXgKPrnLyebSqQd/abPK6GD2/Xe1DlDOxHYrNyxpGgdWiBhzKKI6psVlbG
Y+0hOs83Bzhz6J59JtD5zNYIh4peAn7y5pZKa/s8LZeHok8FFm1a872EliycoNEVHARNWNFN7OjL
Umb7f1tScWHZpjv5jrB+CNwI6/I/Z14dN7FAET3qPklvNXJ3yGX6JoN/52NMmEcqb3bGE6Uh5Wzu
T6WDZnwlbPhAsBxMLmLVGnuD8GvrsHPPkwuUjzdqQqSJ5fUP8JPARycb0qLffbpYmf5laezZr0JQ
0vfpcgj7FrDj0VPcPfbjdrhYkFQudF1PcIsf5lI8ZeTUrwl/VulqhijVBqAVeYYIKUWbJkeKkK17
OHk1fPfTKLML3I5g7wrxeJaKWOSFjrVlwNVzEGS7Pk4CbeNMHnS9ysQeTKzRpd241Vz/fC6stmCe
vnZgm0YTT3G75g8m0qPIyuYgc1ZGYzlD6VR2VSe0Ul1vIh8x5/UraqfWAKECir4p3Qm+bPN47acL
R3tBI004opS0lG1g1hboshP+41aop/mR6yYSfAcwAjEO2ZUA0fcKo7Tx67W3+YpB4lCcxyxYAhLC
LAuk7amyhEV/TNB9TlUH0vuOZSE5rophKb2JWv2Duwvzmzj0W4ECsxlOngdizw8ZOwdOCIw4XHh6
TNP0mCwtfERMUMtGc2VYKqcPpB4/M0Btc07HoSjewnqLy3pkIsE5EVekXpKx4hu1V1TcUumlHfDD
a5hvcgpecH219GonVK3A4fkeDr+e+a6EFX9CI6kAzQCYsQkbqjj1krJWQ7wjlm02c5wrPZXoPiF/
sUCINga3aYcg6OclXcF9DQXsbW2FjwOW0rTHGV2bu/jXNUHqNZ4D3feVVmuMXIceNi2pQOdMf5q8
RlXBCTIMVcHotD4jEuSMmkpVk6MmERXdNeEjRCxjugqGmgdqScqFonpPrhFCv3BV4OM9Zu9FYu1v
asbwX5PwilIUMfBZ/SsqAFxugLkGef296YQaDwzLsDuh/b4WLNccm4eGJ5Jke+xJnSilgB3B6ZhM
kuotjUg+pasL5G1rewZQjUajgi0t4iZmlbBT1T9jrhZ7+J5Sfp9yHhske+P+HvIxrd0e1/FRp7kH
da6Ku8B+edkVM4z2CNrhqf1AImeVOypZc2FUGozsKuwS13DSDhpIZDAtIA0hJVVSNTCP4Lp93h2k
xdH2yX5o3KSV+pAApiD8FbsdURDGnZ5r+p8tWl6zVD7D0MPZuy4fv+ozfxCxDJTUvbbptmU94dOe
iVY1NbNZBLERxUGmyaNvhD+/H5q40RjEhp07vmDqLRnC7DRKCTY+q0ahByZlHZF0P62WdArYlVAM
0c6K85x4485qLBPCV7A3cim3OkfnHquQ04JpORZeHJ9zZfTP4Tf7lC4B8niNv7o7Q7SEQP9LJdLf
X70sFe4hsOPaKWkwAO8sb+d828szIZhqCdiQZ+5CpzZ7QaqoozSJV44gv46F1b1a3grM/xvPfXXx
N1NDemXZ3GYyDNNPmcuDmYWNXYvYiMVE1fqBy0z/S0OAj7qYVVwCoAtjEB5vYKQt2T4tUSpba6RJ
kGsOjq2FGtVwzPlnUoLKfZ1NuLGAXuvrT16UczYBn7k5R7CNmgUTTkrLZskOBm8DML2gw9koMXba
6h6pN8ZEXq6LjXWxTzfkZEI5DTSQbQtRbgdL43etMTd8GRY3cm/4eWwHrOnSFrV7C3Nu4SZ/Yu2F
GYJdnkWyrC6kEe1On/IypQZup3PNxiOHTR0+pLYdwWFuzhhFa8DWkqldLsFZQLK0gB1BeGp2NP6S
wDxJ7V/VzzUjy06aFv5M7nI16RGp4XtWfswG3oHOa3Y2uyofn3ExDi5FUIjJckB+/z3Tq2PJGlcs
0nnhYgujq5sfYeN85APtnMvuSDth+3UARbTzifEvb4wZzGj7VFbRZ/3/UN5uYaN+tfZxjzgAyL/d
z3b6xqj/dmguaLO1oFIHs3DCzaIKq85UfBJahdgegMON1rxPM/CzrpGnVDWyTTaV02hukIUJloxN
UYgK9fyftdDudRte3xPh8oErbdb1ke+SQu8AqE9aWhrN/SCZoQ73vY7061UNRljLvgfLfh57G4Mr
M1oU4T7XGrOZeYS3hj3zDaSqUXy1dF4CnY2G+Dj5hhZ/mFEX/WstriOy2WTssagRAMlbH4o7p4Xn
VBo/zJ18VlorkG1f8qX4gLRYdVIEkUFLjMeP2WzdJ4th9suIru5GuHlGkKUbjvZo9VzJmLg4yo9q
wom8xu2whqe//TTRYTQMtPXxmnMfrnpSjPvbjTKFjAZEs6BiMihqi9639NjaIFQ2VHccg8biikCF
2ipgKcznQ820JzAdhz/ut0ArSDVYJCSWp8fQMg2EK+Yvm7kxVvgqDZPIKQZk3aajqfX7Q9sCL87Z
DvQcsZGikU+UUCPtM1LuAaaXtGGm46nL03ykmdsxxUHLRAzS7rcrG3ZVbMtSUNkKLkXpB/GRtTn2
bKRrZ9JgotxCzPWElFhVbyP9WFpUiVp7Sl3g7kE2d0NAzQsIBSB7q2DX5Oviy0CnL9J4lA812Tbq
70OJlAcNwS1tithXbJ2vLqjJxfJBb1dNd3il/Pf2Iq1QZpQxdXS8MsJ71xUMrQJIGD6q2qy6j6iw
pdFzEAgVM8S5KcLuQbpX5Twlwf0bxgcueS1EPMxsmQq1AkO/FSDn0Cd8kQoWKtxEq09ji7P7vOYI
DsX+GDW3ioqZhM5m4RM4ei3NrxwdCJoJLou/l+ngmKJsW2jU+LPRkf4mqdbYmd7C01hBpmYwX6QJ
STCBCqt/otFpyS+xO+yVM3EjxBF+lo4x8ocfjPgntA/sbA53bwM9OvLaS5w6/wfg2WmQ+L2ySc81
6c2EjNYvIQ1eDUBT5us9aBj7Fo5GL+HzuvL988bT5R0Gs0r5kr+68r7FYuZLMIXN2JxHO00gjTk7
d+PzKhew2OFcWBErlhnT16BmCZBKUkeJT3AkNAOTpM1anB7U6zSQvWNUhQYEpSAGFGfoQaShJwjk
Ym5EIpoeX637kn+QEDE/uBHjCD6GwUkmSoO0qL1wey8bGMP7YZUaZefGylZzWqI9jmgUJ3qej9qi
n+wHgfhYV7WMV3jrBjzBY4u3F2yVQRDBXcO0mAOacMUge3aCAzvuUE363gXUjQ9glOk43d9OEtsx
nDc+vpKdbArVSaoqY7WlG3kmqvfFvfkeZBuEW5nEXWr595E23tnwOuf8IwS55gL4KoFyBqQ2n+tG
h4Sy4/sTY/PmwC4rYwwR590kpbk6ZlfZLfzcSWOuIGK/ZWqpySyTcGUYi5rUZJjmt+mPnSCALxDE
vfyVxc/voR54IOTAzD2L4EhODvk/t/bTbodnVgObjJBeepvtNahppTITUuLA8UmVTbme2mvE1j+4
udnzLM0iJESAt2sqkezeK8XHVhh1Vlgzy6aoslVqzAY8LJw2jQO5rCoUuirWET6pSCB9y//0NvB/
+WraJzoBhOKKk2571f9Z6AzjvRPOCK8VQbjv25xm3z2Jx93i0ZlrP1sEeVfw+mezwcmpC/1UxPjd
zoKnag7AGGC0Wr5KBGY9X53FC5zqlx1MjgVKIB6GtdCNXu4PAJndCU8aLr6TqAXhC2kGVll+m94t
uXriBAOODX4zSwFd5IOBF7O0ddvWOZsGPPk9Xfnt5NGWtQMn2wre9OQY2ixb9YRB0TXmj5m1Gh58
DlJZkoz1fH25Ojno+46lSXPnJ+tm+4Y2V1DNZmzgPAlK8gnq1zHVgIe0ve+rg9qyIOJjtEa6XBde
sDQ1C7IusWBYo2I0Gu8MP9WhDtD3CDsoKK6oKW7fXDJcObfbspkcxfOMkX3/EeaVznKcIHgay/Kk
rqWEM4YPonEvnJIu09vj9t33Vh2pAwYXI50SviKSb9UyJ8PkZA8ZRc1LykfCJdX3uNzHKNnZF22G
VZsQL9BBrJPwkv9AATr5NUL+57qPFzcF9llBGOuQ5Ng3JNcW3vxyy53SEc+9I7K8bOnlKAi2vBu9
6+iNec8nU8WCkflSNVleGqLeQyX8w7spjrOTbmMZlV8LBBrm06vvD9dseYYVj0fuKds2aavXxLsr
rEGH3scWvv6nV6Gr20Z27hTzJOtavKjsMcNTlY/NnWXz9wJm47tXT9Jicii+WifJ4tzVUbdU6NJ2
6WXb3EeKITVVoSYERmDuY251R+bzYhZral9Ns4eADRoTpmR5J3KF9bQMnat7UKPjQI2juaiqRfYh
cYGv0enzt5rphrQk0aotBn6QTASMOMrBCG1IFpMZCaXjJuAGJgMsxNuLIF6PfFPTWhSzL2wniDXM
Uaqq1Soz5U2uMZ00kwYvKmtcerVZvcBbXQEbTZzlh1whnS5mRsrh8NUC1bY4u7CZ1DYUVjLqClzM
YKTzEsASdjleHeG5NysFWiVaHK9O674Pkg+xoImXG1NFd0Fg23Dv9aCGdhMzjbP546Hzh5E85r3+
Pfe5dhRJbkYLX5f5glP9/cMmskcktfMVZZTk79rWUMS3sKdnCWQQGTwNszsTXaN93rY+0+0V/swV
MBX+byYUIDT7jXYe99AFqkj8kkqnipNDe6QHqrkarve91MymMhY5C8gmjVc+SI51iTV0Gf2Od0Zy
ocSApnkjPpd5Vg5A4Sgn/C0+lTdbxP2+IumfoD/No88q2NefCYAZ68F1u5LJZiKR+V2D/r1Y3dHp
zCqrLPVd0L9HcEkTvYYXJ2RhBlAL6zuXEc3DDRaXmnWoJKbndzfYSlGcO+OdxPotv6zi4jITEDgU
PCytH2l9Gj8fSjZfJnJRfEa5fuO+LmyKGnO/2Nw8vx3jirwxlR7Wrce18Xg3tey+G2nWBSg0aG8n
MdW8gEEojq1v4cNCrG5prFKQikP7JBKrLl7MzYPsrGUlnxuvAVRPZd8vvbB/xfLU+D9u/AGeMwcr
0UdSguywBBDPBfaE8ReP5KTnZ63JVSYpOdCJ7MTPM7Nu7M1sBag1zNTImq/88EnTqK21RnZ4ldTA
VZjCZUV6qr1zrky2ODcBGd33agyegjRUPplkkeovSActioZT1FVe6aXwwv2Fhat4zlJa4sAI5hQo
Y1BwcO+eYxhEMjNbrfuedxfN5YDrP+5s/5ViWwf2o5Sv2bxxApsjwHNKCllPNjM+xHMFny76wUXA
YOxx3sV/mCfE18XzQj9SO4hXPhtQBmJlPNCm0zBiwhlmp0v8LXEIzFkN1ytFjtaN38MFvOqtXVT9
auVsGCyyYu7YMBAfAhEI0+TWYboEjisc4yuPOjOubeFs5s8tRNqyZJXCs1lh8PMH6ugzH5aE3p0o
rlnD73XHCDL6D/GBPaLqZzMyScp2XIJCcJYcH+d4rU7azir5f8jHrxzDBL4YLb48Fkl22uQrtTBS
B8s6BYo8pvojWL7Un/KD+xIfF7JY43E3j0smKkZbrn/RBe99d52nEcXII+yoWsQYu/3VvdxfgpWY
dOAbcHZC/DQl0PH+I3/Bh/5vpteAXp9aqkmtG9iRQWVK8+RHZQV8MedKLf6q1Ue8HqRTrz3OtZ03
tDrfNhV8r7c4o2MKKrC4zEl5gvK0jvb/qVObnO475tPYFn2vvH/d+yy8Fq90/dg4KZQRq8MLd/DQ
RVRzXenhjdVDHwA6IhnIPiLhOjMP30OCILnfmgHG/QxjXhfUj4lUhRKIgArshp223qM2K+JLESXr
KSlhurTuKLvBcDSIKBslSsDROLd1V55TgoR7koweFJ+IvV9f8X6kxuFNxq7e6d3k+6VaHOj5Fx8o
iOf6hl3S08qQ5eCo2MYqd73QiGj5nCbANNQCsVY2uLJfffayJbyRMfzr9qJC6hc4QNjcyvwMNtlG
+5TqmsxH/smH704zQTwEreHtqyeXCBaG3mZ3aEJMNlawufLvPHX4Yw4Q+sM+eekhQOTrb4QnFLGP
g0lECnJe8NJXM5kBHt2i20SRMM9Flk7QPKld4RjxsuZaEO6yv4i49WNKwoEjrEvOSuTfW4nw0xM3
q07d0R0xOZ0KR/o7WyAvDht7mroF9RKteqCvJA8QnAbG7EtwsY1uGaCBAzNtjJdnNgqh77CIEJwL
0d0CrVHLJtwvYu38GbDvB7Bey3h/NEf2m6/8Jwb9YxwyPcRPYNUzNNfafPATRxE1lQD/iOCgb/rz
LgQ66NoJQJemIwZWyqYzv9OR+vZaojmXt+JYg3kyNRHIIrcZsr7yD+lAnZt9Pb/APDk2xztnHBQG
LCPzMHkYYJYW0zmfCrGUQukioVo+aV1SN2YrTioBt4DgIdXPr656S4OmAZf1nsLTZdwli2II5Njo
FdWvSH5YP4HetMYobKqEsxBEH9+bBWFaGPoOjqOi+4ne7a2LxDjqLPNiAqA71Fp9+3B138Gafosm
Rux3zSNzhrmbQY+4iTZsv9Pw8CcotVzqP3FtuNtAyffI8pxmVKz52DDZJLD0IUfefI+dDq/GInPk
xxZBE0tWfX7F21iEMUQLdUzuilM3u48Bbo+mKLrrgshRU/1CEd665lLuck/I0fdrPRYqDZveWGS4
ODR/tz2BgBAC50T31CHoDxDMA2tKz0Uab1YgMmREXvnQ85n/JuXhKKgXKBH2CGapwxCRSsG+fzmf
dLG+0vYRlxc05kUF0aOTsUfaf6lhoC2piw+ibeM35JczzQtOxel1WOlD8qvN8uKxmATd/pJ9dPRv
9/dRH3XM9hzevEXZzI1cAxS8val2A3UQEo04gcQszvHk2to1GeeH9wNd+XcmVfiX7mW8aTj2eJYM
6NFtjX5CgueOJowSXuGg2Grw3iCU56ino83XhzPjDP2Uj61xglK0DZjUZkGK/EYJNQNhpomaHSlS
Ni7JbT2+F4fWmhB6hJtPUQEybC7p/aF4nMQReFR/dVGYA2TeH4uuN1seSpcsuE5txfz88/iEaOqU
9cpyQjbdtPGdccnD/8GsPFeqRUAO6wvLCqXMx5b+CHSWLmVPzrEVntVdJywcKRa6nnfsc/ofkPmX
arknf5lT+9V6mJafrV6NUKklyLZp5ROxxoDKqLSFt59/2m4c5E1MxHE6p7I8A/oL58wh1qAaKZFX
eOFhv0CB1ajinSMxZw0eRYddzZibCIE6JBjEXeEvTIX8FUSD/+vzIeqf8W7wSqOQI+msu/Yqh9VU
lIylLgDFAduoeonHqSR4srjZFM0L5Ee+l0XF2BI/LM19mWmRxuOk5Apwc7Jyq1K72SgdqXcevitT
syop5rpyud+nj2ZNMmhWFvdwkRZy0j0JV/pfS7OTmiwRQRQCjuNmwDiFkupY82Ah8pp8wpy8XWhN
aIZY3eqP3K2Hte/QvUH10i+1NLTKJIyxKDOYZVJmam05I/uww7X47oGOZZJsKvju/mSwdNRCgXmF
PevEMvsVSRge1CWw+LmvSXAzigyicOmwhEyMA5P2I7ibQwd3+Pw21UNT2OPTLiQWGuYYSHFBcJJi
V638ardchvOIlIf7iUiecGs6eBPuwtqMh+D1gBHCtlfrbhm+dTAnJ+lEekl45/ygeuwWIQjYGLkq
3EtBjDK8pHrcrUOZKDOiXItD10uRbs7ASP6OMbeRktwFJqIbQn5jUH+mF5SlShkzEEMi7njfN3i5
XWdu4KU0nZCrTFg/xSaq4XcBkZyVdJhNSJ7L8HvTIY4q+gtsNxaVT/5KGu4MiLDBoOlgRk39OQpv
g6CAJuZHqMVlrUbeq6iOygQHc68Watozu9V2t2DW9kohfQtxNGngrEMRhS+1RzZ5YTYSWxmDsIhY
q0LuZu7ZkDzPOv+UVviVRQuocT8Y+YyAnFxnuVGCccP/16P+39sgCkeDN/oRmgVMEZa66qmGayZt
6I/FF7R0kefmUD76SNzZvo/GbTKWhfz6/TmYXD2RqTwA5phFeb/ugQNwr5e0GOv1JMCbTJ0vz/93
HesnvQN7uBFIq8o/B6MGbb8MvPmupSirv4rAYD2AlZYkgncefyAEVHdRlkSwUVuwPHoaI3MzazY1
4S42w5nlJ1I8JhPSTtqowgRKQAGm/G24W7RfkmftbWKCgzXiXLhrD0keGZvPgMizLoDOIHw+T+9Y
/7BiaDaEwATftS4WIh0IAUq7QU3pLFPUI/wUFXG3zy7gmt5ZGptRBnRgDAecjMm3ubFszxM8kfRb
ggmo2JHs/lV8w48w2p9FVuwNABqYzssfkUzxPEoWGZrIl8LRTXVTKAJh8retp27pNMcUMigwJRbg
3zfdRbP+TF5AqHtOABPd5XlpBOtBfYUkx2MClI1g+Q7G7h+Wxe85wCdYqA2rgl0L7BJYZcQc8B/u
WjzHFxVzc1DVG9tdHHrVQUquCn5AZ/dqx2CFYmWEANi/ZO4WMCYU9w98gusD5/J9vLWbBquDsLy+
SNuciEeQchRKW8Gdid+oPA3/x6zzkwcG8Pd2EOnyuNBK2AKyDGSOXxT9qlX8Gz2AZ01km8bh8I4O
u+nmzY22N8rA6DqnhOGXKHFw8nZ0SdMDTyirdDwF3sOYajpeo3OZZcmPyemx6aiafRaLomhjglo5
DsjBBnlowSm8+Zv23+rZKNj7ptbCzXYMKE+jL0zdHXM1LooTjMKhSVEH86CYNS0krbQodgRjsfor
wG5kAu6b6cHtfFYWTXbDiPkisd2E+0qT/TS8BOimwFzX4ZcJ6cuc7F/nLo1czXga5+tqj5TU+1A2
ZbCLlpKAWNBK5kTwQZFuN56OxOiaHkH5mUBk+Z8xy4fbu9HE+rEsp4ltjdry6D5ZZC8jlLuO4K0B
N93mVp6ncYgPYr1cRkxth8D/yF2dPOlg6qdVbG+J/Y1YH6nz4RJJ3Y7PsHCSjkEBRhDQt6SInxT4
w2OGUfDxmTD9+YvUVtIABGjb7G6mPMib2Z0dQp0jmn2LMKuWPhzVYua3qL2qLtiYQK6Zs8VRANuz
eU0SD9BNgh6VMmI7kKBBbC0/wirWmkE9XBQNkXJIVG0ToTvzIWhHMJUrGBOgQEcPNybXf/0hpeJ2
rQPmarc+y5duPSqREIgjfpxnjwI8kfu1XRxA6I+eab6rPHAxo4GnIpIG9BIOI3ctSe+wStxVfdz+
yDAfHbl1oKr7/VvhgwNJiS3OVpuXcVIXxxHB2/yI5sOKZwQE1Mpr2oJwhfVw0wv0YzRyI/ji6XJp
Bm/pIdlHQf+IjGw9wOtUeF763GAkJ++TDjEcTnNhChTB5FMhofhsJ3Pbc6ReJOjjlwLIQd/jz2qD
q6ATQUDu7mLiADB6uyoqK1fSn37x3FOaR2dYInS7Fa1tyc83kQecwfWedFwCExBt6joeM3Ub9n+y
0IweAIidMHREoZD4DldjZDKs0WeCFpSvACRYHrEyCAU6q7lxwhNtp7FsaTkKtZKJxkOa+dt1B+up
wJ2F6sDvSubptzbccntpsLCxaUl7Vvj44/aynRRyb+FB18PiGRMoLDtDIevjvcgkEaPYDKNuoKa6
02Rx4/PhS4La+LOk6IkjbcXRMxmawBZ2pEQ95R22DmkC0RPDY1pZblNQ7K7sycZwCqrZWl8kBxkW
0HlZ8cpdGCD09leIC0OiQXq1RzQqP0fDjEDuHi3rQvnh+/mH/qMzZy8abFuALZdwqtg6/DjldraK
7UQq6vbuj0rHqIHkbxe0yvkFZousH7vz9BBZh5kvzIUtOSl/Uz+ftTdZX+9eDK6s/fRrv6EyfrnM
24oiWZwVUHu9fsxz46FsMW30d2utW8EoGHnR+mWkdDZxJbonLb42KEXihrV/nZCsMaqJZa3/biwC
zR0J8B1UMMSIOkWc4X8pdHFn7532A7kfyshAwLI6vU3tmb+kM1NesPCAW7M9hDLl2O9TinfUbKmx
JZxbW1o73IAGNUY1CCebecXoRDuwbPgtuTvTq0WGmiBCHqRT2t4DaQUsVZNcvQFbBMxfJbUs53QX
Kdg3dFn9joeqCWA50ab4LY9yjNIeZrVzDGHbtUCl7WLVyVziou85nV3lAHEqMdJlC+RUjUJ8yVN/
RgXoaMT/HvFR7MDcQ+L5s9dnq1P96B8CgsgfhluMtMpuok9IfYLuvokpBiAEy/PNnerE1tyusnd3
RBCZhZtDRH5R8lbsFlTN8dKEOKCH/615tnLSlvfcoIMsXAOdt7UE20dVVjG7ykMnYuVVeXcVJrrw
rLkwH/T9kO3pemOBy0+R/3oTIvRv2C+833+SdiTUDckskEV0WFeDPnN4rbsglZsDanOJnXt47P0c
J4fww4RUz1/slyo5TQmiPqYvrMGS+/5IP793S+hcpanhv2LupuZTrWhYOg9G/rSSSFF99kZx+rJr
bySWQHh7DMWrBaVriFkbXgXquMup9QbwRq9cf8fDycyJLimdcyf98UOqJLlr7jfWR311GbZwSzLk
9g4OoGUD3hwW3sruMCjlibSeVHAz5ZA5ZF/sEph1iqtOhNfFiFh9v49pNzMPzsikUttrmHi+kvd8
d8dbzNHAeqhOL2iUWJMdIRu4ZASFlbwlxcRxSP1xPqqVe7fQzKgQetSmh+s+0FdlBEybLyX2M+tw
+DSycbp6mYwrMFq5J//32pzQUMSaZUcI+dHw05fP5bVLvx0OfLAxzD1cVmtUE5AyB/WFkmwXem/B
U7v0IfYMrEQkkjavqawETgFCB4/DBBreiqK1yfLC/6jbknBjh7ihSLKrv/FU+6n0q5RlnulnUOwg
XUz5SKBJmGCrlKtvNQEfROPjGLM0cgA/cjCPtYd4nU1cnzV2hBzLAw7Epg8v0ciMScnejf/6HS2N
JR489GzKL4vNUowqxEsE+1rMBcpIqwccWjvzIxVHye7pmCifc8WIjobDNtlwxzgDv9bPKZO9bsI3
W5Fs4WMmFZ7agU0+tZlR6r6LV56hV7MCADSz5KJRoHWHdk+ri1jwTTSKlnYKi/PcDnX4t4ElUIXo
M1PDgOSoiE3kjrF5lknHSCAAvJSzl+L1BMpm1Dnhqu5NOt8mC07fY+Ld3/wm+lXkAPqo0gnAMi7/
fzexFGiV0aMgLdq+1KOIEBxbvivu+AH36Yr7Y+eho3k1g1JUlVnfmEAdl3phUUm21HYsVxujvBsi
YCsnUN1nLi3RXt0veLnIwEHsfoC1Fl5xtSWbs9OUIyO+8bM1x02NpFsLcxqYFAd71i5NwRBS8jlL
lNG+4ubszCSSSoNqJPxX9NkI8dYvYMx6yaGv2GS6OWkVZfj2qbRnlIr7TeGW1NjYPzkB6G6R8Ewy
O7zWf8qLj5TU+He1uIeKfrRW7bfoXKZ6W+Kn6bRwGwCIxTWSmFacVMcj5E4L06cuHfOF1D3wQ55J
tLZZ6Q/ypx/nA9x1kYhH9IMbSxUOHoSLsFy0jr+7o4W9LwpGwIupc8z4jK1qyIxZl0UwkWqOqrZn
cWQvAHY/o/rbx6gekbmUbiLWBdRCIOrgJ1hXXeYHs2G0Cnppsi/BJTAYoSYNhc4pZGEw4FcR25kN
el32Hqlf3XTO/7QvZBK9nXdEN2a/nG09iWA1fdYVyGN67q11gujh3JOqtbrPD1Mc4aRK+76cqVOl
KJOOVPOdVz3CcA3pgIDX+uyKTnXdgNcw4em+TDmcEaOeNNCgKWEhBWChLADDUbgmepFf/3L0Wwrn
XJrUciFhE9Udpro8WQNYrdcKEcoQswE0NJALIM8pQZvrnWTX6Zk35v0wzSbk0vODTeMZcre1oxWV
8IvDZsQsMoVXZdjHfwHtzQHLqH7szVRPFSNwNQYinSWPfRTqcxOVCmxpJA9PyH+rhGuvvLaQkzlN
hbVMANPXqj/dvHEVXXfSuQblBycWkLYvZaDK+fKNk5Zx9xiKYKFkAbkgVfhjWV+ZS/W3Bxg7/bi6
dQEMb1NY9PqKkB4LH2CDBi8d5CfbGqWezf+xITZtR3qzBvWdYBvLd3HurpbHwO//pdf0+kmleFc0
RIoizCS8MqIlBSV2OJ0zN7lfW9A46ULT7WIVud+mu/eeZ0ClK5hKRKvXfLSKThRbkg5QaJE7PHdF
Fmh2/HMwTe8Li7ipM5bX2wOca7hVBKnf6aD9mcJff2GAdobB0iR/9yJxUWAx5wb17A5oXkz23+2x
hu/ilv0cA62lvLPbFsDQlO0xsmimpVdXsLcGbz6eRY1O/cuqFS/tggOhdGM1wCBZPdjhvuUuK/qH
NJsvkyr0jbjBf2pE92K5ZQ3w4OhzQtFDCVHMNkIq5oJNpaMavJ6mnlaLD98cB8/AxC8sH5AAsdCw
/H+qrIpCxy5GrcT8hIE34tkWu0SyD8+NMfi+PYkzAsSHG0gSsbx+Gix0g08QejatMdrnfEDS2ait
hCI3sFTmF6ApvNCHrlocwNcXkQcNFEG+hMtfoXBIvqC4URQrP3sJpnlrCktBK1xhhmW6KBbVtqPD
sN9LPIB9CtcynY/NO8doTFhYV+IFGnoIi5zeo9HihEampd89SlamgKJg97D14ufo+ElERwLYxj8q
pAekYvxIDls4AX0n/JJ9gQqbTbQdmtkQxY3Zc4RZGUn9KTRcC6XX5JbHeU5/CCyvzzwNtD3q4ekL
qQ4HtpOM7PwWLHfbxrJxYFiXDgt7fAVe1lvwcc85uSKe311ti0rl8J5c7KEi0yQaH/6G/4rZrOO1
+c9pn00kxFcUO9wv/+Cf18gLdGAc4pScy7h9GquPUNAVmLYLAuzu6cAbB7Hol7K2Q8KIw4JI+xmZ
iF34MoJWlvzwpYZ4VFUxo1iVnOeMjjXaB0wAw18Q6y47ww2YE9AjMJStkZpp3T6BMPniiMyWuiBZ
HQU1Sc+aM/0ZW00xCMSf3VkWDsFjYUiJnFAD8YiCt345TiJ+TdPTb5Uh9Qt8oJQ/e+FrDX5HxRu7
MDETQHubU2FzT3dDuMqu+RjR4ZXlizKP44RLrkvnTYByYuJcYPax9EtyGO+neyOGW+lDE0zXYizR
SoAp72qQXSD0Ma3EBcchgg034TO7VMERYNo/th2uj1+nObgXP0CrYHwQG8SrFbj1ho0KU6DChk7+
a9UjX87Fd8DdhRxZrVv4jdqtffPcq33zD82G6M/uNNOzrpbKWTG4zu2hoC5G+Gt/CtA4191zo6ri
vi8w7iRkWAYhf4G4lQg0V4zNJd8bBm+QMqcogEePu2BCa4AOhPEe6HY4DNvm4Hb6E+WDHs6b9jnv
s6lOqawhkyuusXmTHKBa6zjO02dZuUDdg6iQVJ01GZt3TNxW0pwi/vt4cJOdKAkHtFN3fRkEBexn
Du+h8Gww9xLx/7DqM8tVyStzHrom4XdEhcvPIp1Lwki9zDEzoL9rxH1tkjsW+Q2Y3Nn0GJBH9yqW
FGnOsq93WBo2H/MivqzDjN8q+o61Yvp1HuhF/3tzQrmvc+i/CATIOMGLfBeHZT6USAYdWq8RZw1J
MB8+hd0J5hxyV0dDiKiSQN0ALmBrzATDBZeBWjwS5IhBTUobkSsWSfFX+/5I/xsIxoXWi0icti99
CpaKNQJ5OvKL4wCFDdDXwZ1irCGvFVmCCnrKln4NEvSpOUwRS0vBfCulE9oIR2yWNrcyJitYGRhu
kxm7StNLyQGudIpUVMX8kcRnYnU3USQKzUP1Yz2RfJDJi8k5FbLLkiBliG/TIBvYR9CDKCjsij4s
KSALHQC619WLuwgjPZRNwxrPRB/kC7q8GimoUxLZKOXgHre39Riut/JSsW1LFTHN2a06YMRGS73/
pAmsA9MnG1e9ocwMzkfJQXG3tcJ6WmWQN1eWQQgHezh8HA3W4+hpMK6Hz+59mDhMjWnasE6nwcrf
IcszOsf/CSXOYRW+PvegSFKB7QV2H3pyeEPV46I87VCpeCQRTaUsnI0/K2KFuujOHRLr1h2uBpZ0
3dZ6vLnhwLnK45mq+UpbtBWpIrsOU8nl3i9GdYgpO6lrmwXjxyzvc9ZVgGyBYo/WMQWcgbV4uwo+
x/XBLxrjfjxAsS422bHlWSRbohhfKHI27sFjFXXhBjdzi2D2kSfwhFBiffNHaYlm1a1nvRugIUpq
Bt80/Ofwl2srn2nUJfJMK8xoRsjeZvmtMKGUK7fVcWEDWFpxQfMnDEIWqodxCHeOTbK+EE+cogKs
ql+avyS3OFwubA9DQ8JusQXHLnGZiQFvrT7UH6Do1udkNQwgI3bZkL4qlRCBskQrL2oLvF0wDE1a
KC1xcCELH0wCX7ikUhIIPN6npPSS6bdTb8tvLEIK7NYA5ojb5iG+/xLK7RXgO5keOhb9J/AGv/1E
3NYrnSN0r+f15AO/kmQbJqmeMtQPfUajrXbvqai9IPJPrBxXmeohDyJmKoktV0Q4ipltt9qrbao4
5sfn2Gf6aJmt9ecBLqoeKu9jVDJZS+q5kRbVPJdbGFqzl1Byx9WEON9dtARsmhskU/UHftqgMyjD
R2LQQVg2u5cAnxqrcEqR032EQmyVPXNHyaHVIXs2QK+Eu/KlbKHQS1KGYa+fmeMC9SuizRy67e8b
5quDBXO/ah7r0jAyIXZ/A5XQAcXxghXFUeHPBYhGiUBNfFc1KonQbICzQDazksYhUPCFHDkIp2Nl
voak8pKbTG2BfQD06avSSNif5qSbPH5VD9tFLApqqSSAwgXhXqevXfIIqM5naAWbCuhOZ/zEqBNj
O+8SBUYj6OPCVyP7viNexi4/mAEFoWvq+Jg/hd2wTNEFt9Rp4h2ZYJUS4QKV+7MW082h+04qSWVk
yyIZxp3mvrc7Bj46NaMicXwKORp7l3OjCcFzsSuHQPuR9mZL4X3rZZKHBvImVDEQx07ULo7UkyVy
SpZO3rAKdsyTlwmUce0gKqBn02f3z4POaMDb5fBloOiW/IA688akDjX/XutXVCaOq79s4o/p2n04
GhYEU28rNHKqDCiN/r8mVvrTza2/i/KiXTqXpdT997qJQTGh5/rjHEUaMBDLYjbihwQtzImny8Ec
WmVsW/JKRAwDBT8wpZwzKj2OpR1PF5ounx5EbAJ0qu0RAAsxYNfp7ZOXdxOI4YYdajA/bpn+rzTJ
Ac6EoU7M2nCpszfYtWFUAPqUt0zXvBFM8iXuSVvlasK6nKSkH+WFnL5SRgnuiN4F+oiNQXzakq+d
8yldNxhRq1JuGFqkO3cDbsQkGbjjZ+VCS2pUII9A8WRiw5V8+k4Ig8pGqKcBaVnzrAh2YOEpsiKM
MzZlf67h5n699LZLTmuvLN+gyaxmRY/g5iwmB2kI/LO0/kquAdrF3iooFwLGZozL+qtHTiyvR7Ve
iQ6bT0c5mVsGNRq5PNQw228Bn6BOQBA4n3lgOBB4jeebXVyMQEkFQZ2eQE/o3LTw1amnTeP7xz7G
S2F3s3qPNM7W/LdtIh5heDAUHta1uLfzgfTne590Zzh97Ai5xN0T9gOsGs0wQegNNMkysUu3yxa+
4MQLhUGfhPZB2KFycNsF9LGy3NKpxXDSZFPulAZKvlGhY2mCL4j+HdZV0vAbQANfjmTWJMVjjsEG
G5refSZkjRxLYOecA53eP3pff08eoSTf67ajlj0K2OzClfjpFlmbXI4/fhgWKSHO5IhyZmQc0I9v
FRQBsB8TP/wYh6TYNivQQOiNqrApt+p+twCBY8/yMn03BaeBNMInzOn3t7QWvVfnl8W91fX3Rc3u
loYlzZs6FtyjPs6q12FrQLJ4TdiJZBFrao4rIN92v9sQmsBirQgN6Cr5mWAlw+cSXenle8J797Cp
4RfNlGWVPeDq3pxqyO082KkZ9yQtY+pH14NwY0xpa2rSL9vaIBMg3BmY5s+QptsgRz7T5gpPFKtQ
64e2Wnxj0iqZuf6d9yu9XEaji9iXD8Sb8UHjghLrfuZ0ebL/pfmOpUBDffzvBXmoJzmCPmbhFekv
Ev/AQbYbkJCww8U1i9vKd3VP2KCUIgJwbrKkAJFfCqIIZ8F/0rD/thM1vewl5+s0mhu5CbKmGkFv
FmTK+QmxtCpCSbXf7ixtKcb4ZYJLv9jvDVV4OHx35D8lFcNoZdUBQw2Wr5RV79pR6X0uXILrB3f6
XXTjgiN7x8hxOY+cx/cqM9Jvz8T1n7YW+8jMa4amtcZn/Ui8vEfAwRE9n6Bix93YakDrhmVzdxeo
f2dtZe/xHvn1kxtiEXZSTeC7pXGctP5bE+B3bpij/9VUdWqsoOhIoD/KbavSbvKJonSQIzDg7QMz
xpwvU87LMY8TbVIbbJvyl5PQgaMki5IFT7BpKONaZl54KfGVjAeLsU3MXZZccR4UziPzfE7Kc3lB
DTENxBbbJbgp0EkJ4C1NaPuAsnO5Cs8ya6gN46dVVwJeDRiorhRN8OF//7r7/8tdxMXize4SICvv
jI2DaMRE2hI3POxMdwQ8dGQMPT0Tg3kk+QqGmqzYxCq8uwHujtSWwfoZsZrSYhqI6+HzvAhpyl/l
uby2n1jkqg9NvB8N/5LWuoF5BN3QRK4s1gX5BL3aFvDPltMEN/nlSwSPr5nVWElsisNQhZjVXxIb
UAdW0YK86Q/tV/+Y89Q+MdI3ofgkWiNZZPh3EXRPcCygUZuQOTQOdWxktU/Vc4c=
`pragma protect end_protected
