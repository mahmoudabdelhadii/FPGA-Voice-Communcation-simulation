-- (C) 2001-2016 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
kOE0iIMi2gxfbLGjHkUO67gZsR7XTtXAxefZyfYOEWPZBaZwznDENp2WleAqISdllgNz3UoqEo5Y
MEewfdYnhuZPxzprH0dVUJIJEN0S1il/eTzgSNepnomEnHiYED4Nmso8VEsJxOt8TwMr3N3dVr5s
FX5GFeaKzNDTuBYpZAO4h+IpWOjCapikAQ8tFLCWy0MhheVZkx7biaoyWyJuQuf9Jpv62uAMiBfO
SfDnRmj6BBSFC646/PLkWju+6V+8y2NQ+cE2pKuSFSGg07l7FeJlBjGQRrHYxhkFxU1QKc0oImOs
Al0GZg6oE283K3W3gg6pt1SNJoIwGJFDFSBOtA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 11616)
`protect data_block
3o27Q2St4vF7Hs64Wuk+sbfRSG9DE669qyN1RDvF+ixiCc13yR1HYwsRIcJg9BmieYoA6cbjU++W
M/jLfuAj6DJqxRKLuYn41OFJpwJH6YXlL4sJs/2TD8gOlRuyE4gXluEmX0PbE/ajJGUXOJQ8M2v/
d2bQRLNQzSxaob7DWwZuVsadljqo/h0toqZX43kTZ2gCC3RLRhBdUw8zfKBFdR9/X4DgCaDTByd+
MCVD2fIUxN5cs1MgaTTp9XkD/LMFR4GjQNny5Hpa8/HODxZz/TDFWxPEH02dkeQJhGXRtcjh7Ajw
MGHO5O9n1R36pYfe74R73Bv3vUhLtULdgqH07P3WkTwVMMpEkygplKOsL1TzqZINspKlDo7gj0V2
mvxYRYd1jH8P22BGjihzcvw6LW2Jmfha3OpBPa6x4C7mWrWG2y1svgq9+ddgvbq9FXs4MsKL9l23
Rj61EAxH3Y8dtwqgmMRp8V6kouJ31YT4xNwHFZoDXYI3siRagb33Ujv+wFejtV5efm7yUAQ2FhHH
aDTexU3G2PiC37/K6SMs94Cko3w5uewW5KxdkXk1E0bafsOXXbVjzxr+zqrxVewGglMk7ZFaRv8y
oRztEHr9YKFyThVQj5XeO/O90Xb1S6sucxuUjt4pZhhDIu6w4Nfb6PmuSQggIQs7MbaMe/5ePXKQ
oUqKcPeTnGr30inC3bQxrYjIEwXlEob/E1ZO6zeQAk5F7l4oT2uH+f81XZR4RWgomPBuvsyMFMPp
qzvaEo3PxLrXQlf4UNdf63yR/8Bc7kujav0Ua/LwuVOieFZtbj/cnoirjZpKVdBXr6/E3OZAO+24
cyBEnNk3BqtCtwiGIIKqreQR55SiLriXa1pXMKVWqLZEknJ7j+nQ4hOOPIjfYj8A5zt2d17BOt1/
PcaEHnq0p5PTl2IQIYYYlH4R36DBk3Gqd3Z2gwZW61a0CbVQctNizXWdCgEWprJPE092TbkFRp67
ik74zXqrJ2Idd6OvrjfVTFdGIoKJelXyGEFDoB1o7sv/e5CyZLd4SHaIh5FixDhp+ZgYJ5cLOw+X
Jd9gIKWrxhZnE/XB0e4siL9zi5FEDz0hRd2T5UlYIYyQJNK5UUllR4T4VNQiklXvKxKboCNQUaPO
/+RnN1txCB5OjCGzeeRDq79nVjLmDhRq1RaQY4qnZu+7IbP5hYDX7yiKRkbZhaiVy8FpLAIItkib
uQFDzB/vBA9t+p0KQCYuP0u9unfqmbo67DQ67ZDl+FjqCNnEVyj/cOGDWkYPERflDwtRfSsWkWyJ
cHxMgK0oyRiDxE5PRaBHOxzBVTqT0Ckpa9zUHGj06roO9Hwef1VDh98bpeOstyqyffF4gF7+tHGn
q6zu7teuxhrZ7vqB3CB48XkrILYiunr0JkSQGA8zHFUBPid01DVMRRahcX5AXlKa+TI+ayXiAYV2
h1uSBzJ74Ccz9WYU/oNmZRc+3zfPLaaNJM4h0bkQHkvRsaUesVmwJnmL/3u6finJcligbGRAWk6p
ZPSdypP+qS6hVJs8xXlZmlHX3JQ6W3AlDEzTHs+TuP45+Xj9XHT8/Yq5ORybFxPdBA3b6MeGnZC2
AHMMqbodnDxAecxjhc6WCq+130ClyH7+sDey2YGMukFpGsBiZUtvXS6HKLMMa5i1ciMLWN0wDUZ4
t7fikaZyee2EEbpdERwgMlZ+zcWqQum5ONlcoVXrJKREBgLrcHAh/o0YXXBbCGYEO3C2E+uz6ZlG
ReqC98m2QNWjyCspD2lO60LHBn/OHxcbQJgNKzEZE1RUqmQreT2AHe/kLqBJZ/tStKM86PqDsd1+
w/7R5vcxOmlXwOtERPPg22SIdJys9Tc2yCyOcKZONMl9aXAhHUvxwsv2nL/ZsXlF+zcJH27CK4mO
GN4CBxF4ABo/T1WNWQeldoNjpeN9FLGugeDhLW3I4k5HXJCZXYiuKfIkQOFw1NM2oCr3ffAewncW
bwlxUgzQCXg8sIJ8+wCM+mbW0CqHvPMEOESz6Pj68Y1Ctevl85CGdl5WMYGnH+csGBHQCDcnhvt/
T4NuoPCQlf4N1pz03vWLcrJBTQfR3FhGkAoU3thNu9yp2VkOaX0n7A69mZ/Y8O9BxuNTABbk0SS7
q+7nkxnRuL6u5Vu6G74EAs/o2Xs9L/NQVIFyUL35ZiEUZmNT7Q62zBsIoOG8HKLRegxqQC7T96F5
9lsw9lZvyzCuBKRSbB8Snn2+Ihkt0/WkxAm/dXhu2vstMi7POY39HqsznZXCKF1KKUQcKzbDrnEd
Jegiw206xdf5oKEW0EQKRjxuCviaiXAJu9UvIZGg6u4edKFzTtxq7ai+r1jz7TG2LmI3suFzqgbc
t8k40bAEm/bq6nM7gsr+IcIZmrV5jOnlNcQ0n1KIOOBMpCo/u4HOTauNB9co20kJUnygjCD29M7/
f8th3hI0fnLTlMsfLFgQfu8BqbqedrpOiwnWi/+PWm3FGjNV3Uky+k4TNJ9HQh8kQa2lhRKR+dDY
GI9eUS0TOWPTrrYpLuaKRm0xl1GpPnFFhdUDgcIYa0Oq07N2sVHY8y48xjeb2LpTwy5Og8fwbw5r
bSwmzmmzJx4pK7DR/9u4ZupvrcahFRVAjFjABOXfN0SoDZg/plhJw8aGw2oG0vuO6DsNm5MzS445
KYpkx33Opn7+8MAr+ALsfH3Dgyf1twcRBhLowozzvttI0eyPsFsy/M5CNbEILc5UsZ64xhC+qHEw
Ozn+UGwqtZSRBNWufz4In5PJEa+XT7MIhhY8jy/ID6jMYnJ+l/QlztnP2tFVN4hfNWD/96ClFVb4
whhe77Aex2bG1SG9WK22Gmao9n4E2toPPr039HiqBXk4WrQEJLFGI4m4mR4Tro4D3S9TYylZaGWC
WisvPwuaF/bl47Afllhgft6+K+qBd4JkTb5/M0waOlArYtuYfpDqEbvTw26nFHhiJC2uBoGFeT60
wpYKeS6xF2KOi/BPSdnd8Qt4+nG2EyJRADB3YZhcsndC+SIy7vYsKUOruqjuFY3k5BcK1znlDsEg
Eb1SMawvsvLM7m4FqPblQaDvsOZC5G2ygnXh85UoNApGQkfFAWLQ3hrkC7UeAZbVh9PhK6O+O8lT
/10r0tRp6dd40pt5eCPfNFKWAP3WY7t1BPpGB/i72yeVuKV+BuNMJ/Pg1FyrohXw7lYRLgIlrrTA
wnA4yiUpyBQbZm9DXyUFMogAtYJz2S9G5k2cdybiprF50Yc1BIjvIxGjHiPr32G+ifgoj6BCb27C
dOJOkNU4AtytfFGrb7aGiFa7jTZmOEjLU7Vp+8uSK3j6rzSmo0Pv5M0deemRltFJLf6dxsaGJQ0R
83Cgg6bCiF3sow8hS09HVh6b6me/5wSDdyo8Z/wZZp0Si5WtDiZll8miqUi59+NhEr7JF0rHwvE0
PQK2BhX0Bfu8woYOyyoGoaooZ5td2zrb8w4xu47RZiCISE/W3oq7Ub9hFiptfAIm22M+iO4wWAs5
rjGSC4UJtnrEoX0o6cZvss7Bto9q4ZR6lQHpIfiug8s5RqlM3Tv9Bayc7v39+aZ7yJrtyII7fj/v
ONsETL9msqX7E9IyB25XdPAmuhX0yDrUBtd4y9isa6GMvN3R+FomyUO/cshEo287imq+VxEpMpEq
n0g4mHD2iwy0dzYWtb9+uDUyQQdvsMLOwUQ2bP1XFI74X5OEFlw2oMWF+hF7FEduzKsxwr5TR8la
iHszToEZjW6v725dI2Q2P0RlnSFBsARr0EwbLfIshOJk42YPn3BiQPZnT+zEN83JsQ0Upw1K0LiA
pZPw8Krfo66Ri9t3xWBuGuEsEdh/6k+rQOBqA6t/hXpOP1dwJM2fN8sOISmkg3qyf6H8NRWzavII
2Y4l8TFqbhLJXDgVLN7Nlo4TcbZ+l3PQvLMSWHwe410DMAIGyKb4bh1icfD4QB3MrzOiZayQoKer
XwSriW3I19T3AM0wUjpFRu14vckb1m6mTWju9LyKFbk4ZmAPOetVavbt5Fx2+cw5ByD62TZVviRD
zkKQ/1Yh/DTGOxxeY7U06ItzT6PBBPcQ0QD/laQlTV+f8pvacjCbSmlBsD17VvKlRQZkykId4o3k
YT4C18fzgeJPjS2vW1uaq+wKUR324etJmWa+sa216/aNiEne0Aj35aZ/OXFzwOKd3own8cQ1eDtj
wYsuIKTTHxwBdzm9dT/Jjh449kYlElX3nYnVu2WAn9tEDWblNybpRV4+gLVI6zZIyw84xXE8ppWm
33/+gY67AKoYLKoF2yIntsfzOSz8XJpsTtaMlCwhmdaWmLejN5n15j2z18MpaN+MmRkGK4PNG8Nn
ZR/pSy7pcVmmAYL2Wd8KP5Fej2uX1i6o0IH//qMpL1iY8lxMpW0RuxNzWKBsTjda86QHP0mEEBT4
N0kxwlSuUq9MYpQaZs2kmSH6RW8dPlC1fvyI5cTi23umg5gebj6intiXmbvxXSR2QDB6uDOjR+wl
Ywgeib3GmsYXMj6alDI6Pv6cKS/7zO/BzaXGKeo+Z+Br1iO5O7quab+7dzvetq6LpJ66Yv4np2Rk
to2KjPRxbCue6eyc0cjIe3SRIa/6RqizJTatQbNxWr5tuZfIva1+Ee6fddraWcOt5zsqdNuTDagx
41qKh2sK+0N10hUQsVl2DzDZ0US0vt70Idlj/fP42GpCV3Ny540gZPPtPcIbJnpvcQPzHkoMXjDI
8lqGpsDc+rj/gpm7M3ibLXLIjCDe4CW6LQ0Xs6DniKBEdNY5DOxLcUSZk5Wc7DWa7PcqnIWGiIc9
Y1nIIbVPp4YNJRd5aUOcp2Z/UMz9vnSLxgTq12o2WsP9hZM8+LE246GH6xc+vEII1yRrGY+GWc6U
EFfMIWU8FCjbxgiyTTki8R51wIJN9JmQ+tao9CANYc80DIMgqYdIQ882EeTEmAQIKjrztE+Adz+y
+YeakkvNs86nsxHOybLvyYAspSe4m4SJnEGrTGL6pl92izz9zGgDgI88XCl6VEhyIFpIM/e8J924
OlVlNfqMolngejEPt7aTaK2KxzdtRMchQdNGMgmzRbDZ0kJDO4QN9HsQxafd9cNJdFsRvH1dr+27
34qgn13ox8ht/YpCGmRniJTGOM48fA3HDYFX42b1uctRQTXHgVwXPKwqb0YGthyFNBhgvF2q+gl+
VpssO9UoKqT4vZdSauw84E7oJl3vKdphXYuStvUgEZwNt4Tbb+E+BMQhwb7HGSNJ4XiCmfDl5KOE
RNDaSlkh0HHP3Ec1dH9bffDYaJeZnKbjDdh7Kes5Hw3471Vik8J7aHeGLxg5+AbtJ8MlHPdjzZ7u
XvFLSUKrhT5M3nps59UQVQKAh/7z2oqAChL7utkYo4J208Crpndjwufz1qacop5rTexZtjF78uIy
uDp1T5sXlmhfdBH6UQru4nJ4rq9loyvCGj34WNbzw1HvdJDjAqUwXTSQTls7JO7c1+fpdah+ClSR
s944Q/Y9pceub8b4lMKAFY1i0w6JResPfLFLWtOfcxgLfmYI57D+LEyJHNHQETRkhez0P3Vzn4pR
rCeP3GhUp1ylwSMlZZxqvNj60q8Dn9g3dUqOQ/KWx3EFcUuzQ0u3I/YZXkwhu+dv2zQz3/ZZih2Q
J1obAiGqATZSOM9zAumlEX2ZlhKo172wqItUjjIKP9THDdNk4RGJ5mVhQcT4BYlHE28zWZ3J9NEl
tWX+j/RX/KM/QT/Rsy2MlPY3FaiE4i5zlSLTddmcZtK27W57VisdvFgTGW441APWZEdYct9Zu5kW
8H+wGaFQwjtPJvADcXuZjw5CrPgOHZfQczz2/m8MouTMIZHNORX6+jr6iQjRT5hG0hEuUgl/+NC+
q+0j/MuGSjo8hlix6LVyGuKMYxLLWy6lDVP5LOGigcxr9qcdCcaDYaj9SM3VWhs72LoOFRbuTWqz
+UGFk3k65dfnEYC89lR3IuneX2heO4WWBuwT7wiCjC+Q2ANpVZTCos0SkYRfd7ij/t7t1B5ail+A
eeS+RfNOxJ+YKvnVVX5qEgFiSRyMQ2ELdfuMV8BYRwEDiLVqnmCXJNqkAIML5T7lJ6cW7NWu5ntv
LcqECmajRdlvRZaEgMQjiw51gUcqTOOWQdYT5aaqnVfeYfjdU7KyGTwzdvvtsFwkYt8OtUxyzc/C
Yk0fcB2pIp/0vjB3i61ZhnZWlI20WydZ0o8zZuQAnBlyFMIUIMrgfkXWq6nm0a5xFtLMDwsebTes
hTZ4k99D86kLUbm8KrpIwljDoG3JZOjtb8LPKlzm7govBO7p4HdlxjX8SqluuFa3NjjBjg6GDM8J
+3S9eOnwye6zfBnjOg4wzjVsCrYwmbufc/Z4ojMhROCbv04TLY4IL/hFVfQQbjZDfCuxAx1fI2wg
mmfDI6KHQJAh6ax782jIVpQvoKc32PlbrEb9oFdhSjDIrBUxxOJlYoQjivw9BusdKBW09MhOAMXV
/4/cCMwAbyIz7qg2bYJzEdEyAMVRxPgc7kBjbVLp6ImOquQnLM6bokDKntYIPun6rT82XGMtyalO
U+8Du8MWzE44QZKspyme8rtYZlVuCnSWfjSDHsaAc0odWhkLdTM4znaLE8Gz2d20WvHlQCIFI7z1
KdpgZo+k0G5boT44ZJ1trUmy8UwZue0FG5TeKNyIaYSxzFQ+rslOcn0OEyoyI7No1RCCPan3aE7t
cbkuki6p1N9/x+jrAtgaI0ydbJIR7Mj6EWyYMtd/Ys7/czPPRM0SFYSYy2pTKysnGzeLG4cL5d/x
WSsUTocmwm6u3DHWx4Pcw9Ahi1uHpcYZ8ivXB6G4vp2LfON1ItaSMCP8NVxRt+FBMvVBok4scBuJ
b97BQTLMCrBi0a08viNNaAlTncIjHnW0BB5miPjpMnBLIV4tBy4FwcLOPTomhtJCjLL16Wvlp3R1
dVI1I0s/AEKS0ij7cYTVdP/ZwO5VxyTMnSFj4nbSGJMNkFScEyUKLWb6XEboQKSb+dhS1nEI8o9Y
yA6As4cGxTMMJ+78ZShdtVSjXlIlxGQftIPZkhCIio8YnhC5+ZwBvXTfrzeIAUOrgbYhxepy8jv0
o6vKKYJb2hfrrrHK0YWCHO30Q2XDr9BeT5KuH4tOTmsSkvDa79t90Al6uDT77KpUlO5kVdVBp8O/
8aPT8gfAKH6ClZAcZcibcOO2s/d/M7r1qmcUZAgGHCupeKGSwGMNdQj6VOVZWtTInOqaDmGiSupS
6yF6xTbTmM7uKi/mcNwYjl9kGm9QUTzJZGFYDXDddv0k0SvRncwBtOdztvXvUlFKVETAmYsMlEnj
83hdQu7/ILa8ZKS4/zxzpZm1JbIaRoBWaUYyQS1sfievn275hqrc+SAIS6WlXgq+qnfSAgc69+FM
LjwcRFQCKtv25CI7P/0Feo5EPv9cQrN1YwIhSXvYnjQmlU7x6HbsoM9XxUwlrwY2ZzgcvJd9Slny
VBEgixjhtvgHkrka39Do/f2Pm/9GP0CQkdlOY9mE3mQmK+vTHG7qR2jRPkhXxtKH0PhwItGY06sp
s5cTDKpOA62Mto01GhZKW6eGQyTjX5vrRelHapBsCOPeBYDJD87n0ydG/QDv8lYPTJxQZyniJfLX
Yl3tyfYQ7eQBdoyml0VgV3I6xhQCHfP6+4euN2way5vym9/PDaboWVDqmsxlrpLnSYoKxsdNgxm4
NqDLZ4hljjTUl1bUlPb2NukmmqOZ76Qyp7dqb1GULFXmE8y3XocdA7xo7XS99w4IYJiZbmdhzjZj
Xcp7dlNFeA35ajkf1eFt+vDtPlecmbsDyEHoACiJevFVtn623vvnVvGVBsPN20xRdMBSesaHw+W4
nYTwa718coXSxgx/J9eRJrnieney0I6NWrq8pY5Hp8XWRgZtZgNbWwPelmc+LoA97QBnf6lDUema
YLLXD0LwF0ShV+zGqTLomjmStKf8juWFz8DRoaeSkSTKR93+D8ejTzMnhv76YzEqBh1AnUOZMpQC
Y/zDRXfCgoCmy19i/ANZ2RowCZntmw8DI8zpq4brNgQnXPteI4a9/BrdpuyiYYMkzkSIbxGKEdX2
c+bMYerNUYHgtVy4JUr/kRqfddg+dTvGNE1PbfdO8L7RT2O4CA8xUb1CD7V1/L262HyFbh64GVYr
oXZRiGCRPGT+SFaf/nU42Buj3pJTuwIji4Ofh7R+SRBlteUFa+MSk8dkgN9boLi+gnl/A1uAVS25
mqT7l1gnE29kOYR2pHoICj63BMvAAt015BgdC9rvfMhxbZnUAsUMx1YGl9GgdlCDeiVDcgHd+ctK
Kl4BCeEk1Q8QjaXHsN6q/LffSnD2XSHQcFk+kC4WplDAhYnTHxETigBK3s1XaCHmYE8zjEHLbyyw
Q+4I70QtVo3FudYvnQzvoK4oY9cQKeMHOR3pUP6VprbxqKdXDdPHj0zH/rsmM7tEEYzfAYUYObdb
1QEItwa73tt1UzGjBgLr78DcskP+MR8CRhsyweW+3F4hYzEHMb0zgClNUaj+o+VTYjaY8FJd6wdO
3NPkYrnhU4Iy4fZo5nBZV+IrgqaiA/dvWLA5JPHeFyYrdsmgf40K8eoTE6D3vqAldn54/sV4+I6Y
6ilf+mJl07AOA2lnBO4M8Osn2t94NyWsbTeCRzFMSSlYzUXvjt/Y/cTCo+lJfvIvd5II6yC8dAzQ
NKODqcOeC3F9InsGgLEoVTwYwCN2bL1qFh/LiyNXgYGOYPlcwPaGUz16AA/BbEAqvxTNy8Dh8o8q
2rfxji5hdlk0IBNXx0Lfp8K0VxWIrEZIh8stf0cUrJlelylAiazQGWmF3M0s7C2sIGqdR3Xk2GuE
4g/03k7BnlsmG6+OS8O07vqanelfTnehZWC4/wc+/eo46t/Gz0gp3ymCsa2LbJkt2hhTtT9rBbm2
VetBht3YhP5zz5A9VlcjhKGbbEBVF7uyFR0d/NgxGMMdfJdu1hgmXQWutPo3nhFmVfTl5PCuNCF1
kSzcwkuSK8vmEegeGXsLx5w1gKeffn/l7CjlDeQcSDFNkz2rvy8Myo39Btyx0Y6uxq+evuXy8g/n
2HL9yDmFtGLBCNLJ0gAUGDvvloEdelWpaGRakgOaMWe/igWAfSFQ4rohbr+7i8SGfyFJCRZzES+q
OqyDiWZbTw7+GGQfujrzw6QQ6Qw9YhWJdHnh+HOGZU1KxKpr4YUu5CDSz+0qEoNSXOxNG60Zmpk8
6j4W+KGxjedE3wZXnrDNWIDC/GBtBt50ClQqRhwge37S3K5zmPmhqn2AJbvb0PpCuIbT8cgcbdl+
bC+IQ3+Tm0rU5ckFLC/5P88yWCG64xvfTBZSH3dAEbVZ6rs7MBCKaACswD4hPhiMv3u9nMqRr70t
IFd9fvT5GAjH7b7QFKJ7Gf8tlqV/ndO2rvds0uq21cjz8wYuijMZAPYC0ZbFYlZRjdy1mOyqZ+C8
kjbTl240zTbT879lWP+EqmhvcBoDx9mRhj649YedvNG3wKXpe47zSkKyLL9kW3cM89W+6AqRmLLD
8rdiXODs/96W3tya6eoprQ9Y21JimyssI20qulwz4a6bdNGekzGghGpAynU3u0U6xhF9iBav+aDM
CMNEaCxuS0ELw1pBnsqJP6m7+y1ikZR90wLk3bUc0/7dAqPzp0Ega4Bzh6rgtJo+6dhWi/Iuf3ee
viJlJdGzRjLowbDMWnHhIvhqD0tEPqQB1eqd9lVU4x8FVCRpANd2Jgpz10l3fk1zmxnY5R5LfHMc
0L6ZyMOeyv6Nw1zyRxL2c//53VCY9lxrnJ9fR1Ydl6ZTgh6YDpbfGTCsOBUqGYi3GurxFgsbb/mw
SepANndlz/2w69RqKUteCTYzgmCN0SVGF2UoVFQZlXd/8Pj/FPjE9RmU2k3yP9Sqn4H85rfav7b0
1JNx0Tv9pCSiIXLtgPD7f0OBwlnjRwYGJFxxbz+LcRPGuEdFFCC1g0R0d9C49D1mPFyJoM2UUcIG
ocP5DeHjs9vBAAqGW8goMpPWCtGn4cZWJxGUqq7rpcCtChjjOVxBvRsc7fJ4yJb4oOF9xip+z4ti
yQe46Sv5YaWglTVrVPxlVz6sU6y269JqYR+/6i3DjEBRSz263dc17ld0Mw2ZFWUm+1sdnFr69c3f
AtpK0UPmyCgfbLKUJ0qRDofrpPDdnyglaroYdWO49fosApz84KW6snHOvyOgm0SWJo9OVeR9kZcg
xhE4c9Zin0wSXQaxitqo8WSUNm98LiwyKysBLkTOmUHy0WcxzQCY9hMhQJPqcmQSmKXxlPRhuImc
b0Mm0d8K5n+Or+VVi5KRp7uWZdvrXjli2KtDT6jhN9WddbVYAuLwNancwJcMuNOKyEkGYjydJzyD
fvX+iNnbeKfGRotHbExxraHJUiHtvPdejk4J0aNvta15eDmOzr3Tjml8IbdibOTE15l1TG78vlCy
nw71LBT5gFEouu6ysUnZE2F1GT5ftnwB27sFcvUShb/AHpyP+QlkXcXebDr/xe2N9Ouy4d14qmX8
1RbG3PwqmpiuBinaC/YppkcBBpSjAdpbuFWswFBy+LIEk3hsGn6BUTHfj37/qTZjGiu39uy4YIeK
4gDxGCJxpf/8OLe8ScNM1euxR6KCtRib60+Cl43jao4Lk4sOqUfVYUMOV8QXfdvwnnp5ehsCrtuu
52jKxv67h1YjJ1phdjXHUUMGdiTY5v+6RnAVMihBdeZpQxuabfs+m//Bj3wK+KrTNnmK6vKn841A
0yahNa8Nb2Vd/3OrGxPivDblWlLgNK57fkQyfYxPwBX3YB57JYgQhhj1Ci1i05Pki4or5UZfCvW/
+9zpJxx1eJjsVo1VL6/Uahyae3WUCe9+oodRTWdDZSSsFdNoB9wI3bSdCVUZAAghzQyIj+lxxC2B
JkPp5H+q/fMWMifbrEr6DNm0AzBBsjsGgz9uGBmSXCCz5UybhGzgc37lJksoodd5xOzv/bebBYTr
969a40lljYLaeNInwswxEzthDG/pmMAJRPeb3gIzasLU9g7V3zQej3BiHOBh8lmkJ6c/nXHgYnPH
XFJzkti3LqKRBsQeH1wTKHPJoMTG9VblHfDmhmKsqFFwrE7mgZQriVzJsVFfxMd2OuaIr9g/MZzb
oC3iExfmLc5x6IbaOQem7aT2P0Ae/xBkHCXKgkGpC1hG/ESN72CknXuYGBhC4rPFb0ihbJVkP0Fu
4MR+V3roVEqfGCFEVMn4OXKhrGD7wQnBPNrmRvNcmkswatUr8p2kGRSr/4S9aCMmZbjsWWqp34yW
lqC/y5e3aOIaiRjhHG5xIS2hahfid44AjVB9U6nCVCejshFvjLnJ4yxV9biZipyhQH1FAFCzYxNU
HZUKuRT53PwgJ4OKMvLbBS/9lTTRQfuAPfP0nYPRh8/dMfG2g2oRmtYIsVyTgxuoIPr1d4W0fP9Q
d3u6VHiWm+D84XnK9nQOMESp9+5gAlbgNaJqKSS076yuw86xt5ybtwmIgRtiGGmlaJEiVf5xOlHq
+KJytjzXtzHpaaV2iWf47xQufUmNBh3htEpyfCKi6SO9hTYwBksW2nlhH6OlLYUkML/kfjpQ/0nK
KHlDUG0X05bLiDXIX1P6Hw1dOkMqp9R/s2N+buqGPooRTEt87xsfHkMye4Gc7UPhxAdXjQzvjr0A
fDL/rHy5z9IHnafoVI6mGL7XaX0ox8TZ9tjgl2EVR3fsHn7/5FXKjGoLQC2aiDswQ4lwHDEu+25h
OnOkOdL7uGlerE/SHbWgG37pJu2CBLgyHsjF076gzGp63ZdmLGWbGemrNWylGmGMmJqcg1sIXmEC
dOYULi64vRKwxH9qcntA3OMXkW1Hoy9W8eF8hONXexxihmukyzplAoaQZUM4d0XMdXhedXSRHdjA
9XYrQ6o7egt2sCIxBBwuKxNj19LY4FByD+jgjIEU8zM6HdUawGqnoWUDHqU+vCaeaG8m/QLlZYL5
aPfHxyL7lUSj054wF+P0eims5RTtxIOn0UMtNS/u+REFA4cHehBq8dXTEnXOtq8xYPAyEsOiTVyE
f1GyE5Y2Ddg9uVvyXQb4YZfSxLIRJvk7cM8YB1Hk+TOwmCBIbUio4fTJhx4k0jPXLc5Lk1V9xXeL
nPeOmSSp7slsuppxkFmo/PjL4gSjbIuHUahhPy84FBZBDQTnLRnmkPverCB0PInvIizlZAxiDjO9
m164C1645PBGttWuiUygEYxUQ58L4gzmQc3jUQq1J5W2v5D7y64slLpCEcVoR0uvYsUpCeqvufu8
+ums0frgBMQSg0POSDTSuXoRNEd0CUkv7e4rP8boFMssuonANUGyIvWPJ7fULu4SjyuY6LhB2UJo
6HjcUVL31i64gcJT1H5I0oKST12AXbfZkzTzU4BJUER5Mz24SmG16SKtw+DADbkUxfs3uy306Xdy
3aiVFBqOWQrH7FQJMptfsqDnBVV/Is6sn3Hl99y1hwT0zoFplAB8/uI32WzkJ0kCjbKTY5E3MEm4
613dpM174A1yo60b1V2SCD6RRrnFtYE34pnJgvq0zT2X0+3ovkOXVXeY2GfeJZ7N9OF4Yj1hP1Rr
/SJZuu5P2wTGT0en36NXh/cXS0ypAlAaxg9olZeAkF+6pyxT4PAazM5omeD3ceWq2RTxI0aE31iy
x/tg4wj7SVxOLD9scj97H5ZqjZ1BmQUmhNmoUMXchY9diOBhSJhnr+kXmxNvTxL4rh4vm+Uoqk5h
hTWQoqVZ9NdpxKycevlOEc/lpZ/1tPICxeffghVDIkOeTGJLLbIGHEJs1I4h7mjPWdzq0NyHgIth
CsZZC7t++J9JubkUcdMWIhaq6wFqpcNHZ2iTuKnp58cx6im/xjJnJU32kflZxGWUREQr+nxtgaAA
RU4JPRZrc4CBL4vbAyQ+cOK8HApfSg4PM35+nj36y+iyZgmioQa7+NalTW+Ac5tPBYhtKQP8RuD8
Mfq5C6X9C2RkRx9Ki//5CI7fWPpcHfIisC5yDt7Rvm+J8CBgHUdt85Cg8lL2oRvRYOVo2xdhoBJL
avO2vLcTwQPpJNGDq9ndGuOUsGzSGvXyG3aeYTtIeGKLDenZdpim/2Xc4rlq8Fkh856NKs2PRcI3
B+jIePkvPEDgw7OuXV8HdwEMbdIaugBu9kyhu81QOapjSrjOppfr8aAEZHbRl+42skF8oHUL2cxK
KJ4YxWXt/En54rOrbOTZf8mlV/E6elmo2cbYwCXs4Z8ISuMbo74Liv9MQxwVoJ+YA0XcXaJf/gp1
4UEnVUQQIv3zGjF4bmBdEgBlGR38e7+T1A3ySY9WQ5cbZOOLW/V9NNazRjvjjSjA6DwPWYKOMz4r
gplJI3QOoC88SCUb/5VM+R9R/lV3P822gzrwrpK2jD+6cQ8lVPm9RQ2e8ZrDXdptnv+HiUpT/Iub
0n3viYOfhUdlH/GafPMuSDT+9+T5XU+EgL9C8mp8PyhuBJ5BQRVNflh4MdIO9hciI2tlB3jKNskl
/7cj8MPdC4wpVVSeKsQRwXzJQus5vGxiReMiZoxWh6heKRgkAgrqgpT5qjfK11qWTBvB4lP2Wqj2
fVA+T+q/zTXXlBDv3aXTh8VkmpSaAmgLDY4yYQ6Lo/4Ke1AuU4SxG/LnrlxpeLJyw7/Kn1cqOw++
UuaX4pX/6v/fSi0BO4A4rzQGUiez86RGBPS8z/riI+q/vjdmt2nVcYMuYu/UNSyQnUs3YZXj6pmc
KCFRmByZ3JJ8pBzFCm9CGFaJNvG8aEvmB+TnB0rRqUoZ2kHspMl2oVzkEXzIuiMhYlPzuq1i4o0n
lfioLFlPOwCTezM6/oXSUYPfaKCkWLUijsT7WrT+WuZDlL1OfED/o52UQqpmzz7OD/ueuwBPRxr2
v5bpwcHsDfC2XCK+2MI8VzbdItzPV9qj5yEfistyxC+YRoztLsNskHqHnWctXWg/7XvgAKTbai0m
P4aPDKq6uy+CxYy/yfL2W48D6inzcJy1gHEG4UaN2QLlboN4jLJYIDH2CXIFFBRvG9URBS1awZGg
gJ0i1xY/fMpPQdT0J/+n46KMN9erxVT2BpcSzPW+Nenhpm3H8Z7FSb2bvrW1qZJL1gRY+mf/uuny
R0YITetVYFh2qUGWfu9bxNymIG1cKqlDDeavlXfUDH5+ldrGW5H2FVGWf8lhN4gn7O3lI0po2L0D
xPErGfeL4+ApzGw0rbky4dC/EImjPuP5XYgBJeISxzHISr7pF9WXb/MkyXvbb4z3ScbavIBfClHd
WNhO9qKKu47cN/VCJMccECTk4nayN7CMhVeo7ABlfJsIDL+oNx4/wqVjlCQSlXI4u+pl9OtVzqnE
wn8r6aBDN1OKLozL3fn7lJvN4MF1By9Z0WUg3Awnn7h9ebHetc8om/YFN5/htdOZumc50s0ZP4D/
DuZCD8244NmYubyQL3NkMz0m4XS7KozheuLHsZfQywMw0G/6MH3ybFVlmgUKQPZYeJFdZbl6/VOi
Iwti2ZZv+HQRW+PyfRTrwA/J2Vb1CjnhfaVliXPk3I57aokIPVb0U4/MnDkq+mhQpASLYV4h0bJD
UhXOy4gJTR8YS9+b1tH4boRdbqAXSeA4g/rM5TM4fibtqgjxKDBKGh9jz1kSO2QQVETPHNGZNO9M
QbEnIX3RYqfWVImisvJnI0V51moZeS9vpzpB50HqaXkW9VpQMqh1oTKvKejkUx1xQ+ABVxnq43sK
vAHTSCpHWM5s/K0Y+S71c9yLTT4b8xes0QljEEAFsdw8xHbumFvhnxRwSUTTM3smQTwG9OpDcrCC
SdsmqzrhWDxAYBCZEaQMY8fcseoJlsU6w/b8q/HeslJ2nVYXx5Wd5xUVQovuxvenEQaGN8GjMi3y
sRN9EQStg2Djx+goFP5s43tMR3jFDF3eM6q14KOxNCUN/KhiYyfEUIJkltN94ddlbZE7O5bv15jv
QB7IfVH0DK+mbcXb+YWu13H+q1olRIlK/lzvexdUieiBFyB97oeXVL8Fe5N3maIqauah8kiPA/PU
tglagzBwk7//lDEf7To0E+cVU2aR9j5xvXGkCL4mC4Vk202UKKU0dTfeJgz5zhzU3ZO/+UDagQRS
PxPX0stB3BmZmvdbpGHwf/Tlomw9hEDslaxSZYTouLXM4G5q3Lbc7puIHA0P+aU79fQg03mc2T0k
PSmJVrYX2Vo4B2Fa9ZVFrcslLGtH4IBvtnjw1zGFBZ5QOl5H1is52SnWrHe7mpH7LMpV8Z+XUEvF
yzxEmBUVLAFhOzrNb0X/GUk5rJzfsXZotxO3rFikzFEY6+Nfywyy61dYIVf74B9pdx6y62S1Wr2j
OeZC4HzVPUMlLXSNmWFDBlo10kUcFHYVdn8P07c4lN1Z17rXg9ilQXyMjGG1RSMagCCPirZDHb51
BF7fDcVlAkZ5w0BLQXrUEW7Wbgh4pVvbMtMnoh0SYTvGJyxFEgcXh4sElH86bcjQr6HbuuePT1Cs
prLFJVCW698Z8rukWQiFs1NBeN+4X1r05NKumf8G8Iv+Z0TXGK2H5uW7TxmF
`protect end_protected
