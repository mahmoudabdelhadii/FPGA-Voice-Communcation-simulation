��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����N~@#�k�0!����+��=L���0�ԴZ�2�Mc���ZO�����=�����վ�	"cqw��a��TS[��{=:�����K��-�մ�(��k��N�-� 偙O��QZ��~rL'�x[�i,mׇp���O�I43��4d�,�H�����SN��d���3���r��m���̨T�I;uj2Y� Er�*p�Q$Gm���p�V�`�2^���,hz�<p��l�Bxt�5��s��\yq���#�@W���f:m��T�	,*�񞭋����_��㧋l�	�\�:��uGd��PǷ��N�I��_����Tuv� ���us�(H�~�{2H�:Zor�Q	#%�3ˠ!��iS��95�,?�.���/�F�i{#���Tp5����Ҥ0{%���2vpn���X�����@l����3dc�ק�3	�Ed&3�ZN O���z��s�yxӡt��v*}ԫy nj#��lc��m戭k[��5)�A#�����8�!�]�Z�s�M���t��w�!��'ÒE�rv��Ϝ�c@<U��\tq+��&|�&X1)C�����r�A~��B�&�����s�:n{p��͠R�X⺂L^��R����c���f��J^?��ܣR�O 1�rV���:��T�4���AD����˩�F�w��)Dm�O�b,�a���1$��c��7t[i2>�ޔ0,S���󧇳Ϟ�ᒨ�-��}�!6��Jyv�醊�^_�(�H�(y^����o#����X��3-�k\8�M�T�"`R�DF6ȕ� �,5�;Ҭ C�k���1\������k�t־9�}���� ���QHF��"��t�9 ?��{E_�7��!����](�S��0�q��w�9��=�i]�1�GʦȪc�W�XC�|�$��}q�6����zf(����լml�dz������*�eLD�*�,�m�]ہ6����D�Gw� �g���Y,1�?�a�D�p�h�.���cubS8nP�6<����߽.0���ό
Uq+��ilP �[K��8�@�%شˌ]�r���Bw�W|Js}��K��|��`�s� >�c�@���a� ��Qs����?�}���X��nr���o&$bB���o���H>O�Y;�got�y	EF�g���x{^��:��gD�pA���T,髢A(���/OՒ1�k5�t
�U���,�l�w�h�O^{�W��6�|̓*���Im6��Z#�
���@�ԙ��8l[/��U���)0aw(���P] ,��� �Fܑ�e��(�N�k�K�n�̘�V���=�Y��N�����9y��� �p#�w����Z<��q�@�o��0�-۶�����[��Vͣ(�=�D�މ���W=-���ǥX���$��T�7������d��H����kr�����>�ܠ��b����p:@N!bƴ!h��k��N?/��_�={?RB(X��J���&�~$Hh,���4�}#�9��4JU���U�xL|��0t�*&�+��
�'5��u}m���J��]T&�� g>��.�y�f����M��Q=�p= B�j���)��E=l�,�Aq��T\d����6N�q;��,��m~a�i�@zy���!η�r��Ϊ.-��z�m�[�kQ*_��ӻ6޴�
O�k���	Z��<��Q�*`��I�(}�?v`G��]�pL���A�E�s��w�t
�nV�Q�{�;�JREBR7_��Z�F!c��U���JN�+��W�t	��NI*Ŋ��F�|����p�A�,��[&�,sVN�~���~5���Ƌ�
�S�� &q�,da)�V�@�~��0�6^��Tk,�� P��>����`̜��l����U�����t20.]j�)�~�����`	���d`��L��l���NR���Q�^�������]����Ҁ�Lı��������У�,*3��q����k�ި��?^�%n��p|ZN��	�����X4���\*�h!�D"�5�j�k���!�m�L�3�hș��\�EJ�[bIIt6U�Ң���B��>��u��F��)2J5o��Gѽ�*�dɪ�R�DP�e�娋��i�4�����$��8�t1��jl�3�-��l��<��,�8�|��N[�l�@��&��D>�#���)+^B�D^2�۴]�*�R0��(f��4�>�����&�~����He��v8�nN�� с�a�����\���_�ο	N��O�,�{��L��d�=���v5R�����6E�Ec��� U.k7+�n����PVh�M��7|~�zK߫�J��J�r�`/ŒaG�n݄�i?9T�u��"�[��,gp�E��G��w�RHJ���0��c Y�������v+�����zo�k��n`�4�	B���8�7҉�[�@(�v�rU	#����"i\F�W�Z,w���7L�y����޳~���q!�a�a"G��'�4,Cw�9¶I��\[��g����W�r6(y�جygt<+� �]n>U#���+��q��Ѷu��n�4O|� ܥ�b�`�&���DV܀��<q1��u߫�h����S��'%l��GT튼
b��^�x ��ᒋ(Y� �oR�>����9�02��pn��"���PU�
Z��H���)�x�x�0�!���ҞGM���o��z��ES�l�I��eE:����m�7�:���Yn{9 W��s  �F�O�E6Q�ej ��)w|0��z�e���(��]�j��b�7�T3d�@]3Fy|��ہ�ʛ�#�t�}-�f�P��KcO` C�ȅ��&�oچ����f�yg�J������a�K1$t�iT��1�Dy`�
��.���:(X���QC��������U_G�jY���u�x�~���� X���[��px�	��2�C��J4�L�`,�z	ۺ�j��Шd�t(�����`��e�͖�l����՗vk3��K��AP��SLe{��>c�5���r���K�l15�h��˟H,O�0�u��E!�����߶n"*e��jTo�h%������}15�e��}��?!ۜHDb6asr�|Ę�?A�-}�e�������g��d��Ùۗ��5����W��$��x���#h�PO��/r��W���W�em�+A�_H��|VF�~2;8�擼Ts�={��~�2�Y��%��W�\f7�"p��:~��yz�,����v4��4����@,�	#[��ϖ�ś!���6E��J�n�̙Wʵ��0p��mr�KE������%7��#�04=�[@I�{���x�CP�͜r.���!IOB_�:.�w�<B0�C��
�V� ��9��������ʌGAβ���8���-�G�N�������c���g�YB�4���Oh��)��U�֬8%u�Jnh��3��qy�����xzs���	�CyŚ�ai1�0����c��70�>S�|#c78���Y]��*�-�AO���O,��~�/� hi����^�i�T��6�c鵤�:.����è9��cwV��7}�<�������`�V��vL�*c�t�p3�-^B�x���X2���шې,�.��Q��9ȿP��/0�;zq<�9��;s��YƓ�Ɔ�ht�=8�s��e���b/.,�/i�����9���hjVE�#4��c�P���t����s ����5��	@8�����C���^jwto_�@D�cR����c�J�d�A����i��'�t��h��덌����a)}#���Y��.Ko�i����&@�k��M�۬�xd�:, ) �VT�F��<���Dq��ׇ�+��y�PC��߸9isy�d�m}H��Ծ�'�r�D�@�-mG랢�+Le�h�;O޼j�m���0+��I���q�B�� �������+��ޛ����n5���&�֢�ٖ�}I�?n�H��_B�պ����-���p�_�W�a����Sz]���� t��Pi�l�Ýt��ӯ�lt+����/�lHw���X��bܭ�&�e�9|�'����g�m���6��~״����}�n�Àl	��3��?��'��Im����`�΢'f����`�J��k��Y�ԇ�+��q:Yd�t��Q��l��xYڲG�@�)U���z�+# 4����I"������N܀x��ȴɪ��=R�i��� �ßU>�4�*Q; :�f�J�s3�ue�l�K6G�~KpB�[̊���PzF�;&qt�d$��a�M�н{a���VT+M��O%�n F�a�K�8"٣	:���f�L��s�e�`��J7�x>���z�U�W����Q�HF���k�m�>��]�#J�������k1�q������R!sI�5FGE�Oޖ�bRĒ���7m�4@fU�f��_���ƿ�C�	�URK�¯�6GSy�+�r Q�r�c�)�V(q�P����}���jfbc��.9�־�/����f(ډ���u�ĳ9����'���.w�O�<\����6&/:������C��`'��0Ծ����p�N�G�`߉��O{k(���NԚ�ﬧ��q�"3�#��B�#ﳕA���P6D���)@�J�PC���f��Τ�&��p�� �3r~ �1�ڪ�����=󠚴�n�U{�:�{TuOr� H�,ݟ�Զ#�r�����C��+2ӓ�dfc�|I�7����ߗ$���,;0�H9�������r���KS�����]�������%��}�'��_Vٓ�y��M�h=�/�m�  �8�Z]����|��*��s�yJ�{/J�
���Q*��+���Vh�;��Mzr>���N�=צ�0F	�fɏ��#�96��E*������>=%�yXڷn��k!��s ď�Au�#[6kԜ��%U�%�U>��������cTT���8�������vKs ��FϦ5�3& �Q�֝|vmG�Gh���;��-[����`ƽ���*�䜾�2�4NL~b!�	?��(Gp�ս3�%��{_��Z��&�9؆m��r������>� ����[�MO��'��� G���!�]�cnx�+jz|~���@���ncnHØ,>�B��V�I���a��s�=�^�u�C]��� �$^�����d^�����ӯ�W����+~�F�2rA�?�W��*�[njcW�ֺ8���]_���A�VȐ }��P�*�O����_H�I ��S2_�r*����c���^y�uܬ�e����/������%����1\��s	~��?e�?����w�?=��a���X�[�U�'�W�}0zj_]I�#��z��g�d�������ú0���
����	���a�lO2
}�úĭ�O�GV���W��j^�6�s*�{�~Q��;��z_�7<?�Y�1k����U�'���,��]�<�z������6�c����b���֩�%Dӿ
�̕H�����
Ck�۔�l$"}:i�ǗePvT)ݛi!=\Z��Ԟ�v=[{m*S��N�_���l4����Aϒt�'����ֻ����8�
���C)��3g�.�q�9�?q�Da��d�p5%êV$-�<�SF��o�ӫ<i�޵� ��|Ӑɡ=V�Tm
ҠI�������CIAҚ�#�n��e�ɇ����6mF:�6��if�w����Ȑs�/i�u���w�Qf��6�~�L�Y��ŭ�bN������}QKէ�e�7�*)�	��Z�;���OB>�*���:��#6������&DK��,�2�@
��3&�I��'��'�1j4��8���ݲ��b���A�u}e �*��鋡*:.:��򨂔B~ڟ�� M]�P��Ә|�GU���,Y�u���BB��Ctl���'7��vf8.���a��QȪ�0O��6a(���?:'���h=��L+���6Q��1�.�޿��[���w�Z�Y�ڮKd�f|Tdc���o�WL�2�M��eu�l�h��Q����_R�Qj��ѣe؉����(�4��Ds�"��K?���g7��ܚ;��aQ^���h����7�ӕ���Ϭ��)Q��O��ü{�;�!�QdX?�n5��j�ޠԚ�<�!{��_��}Ȼ����{�|lц2�f2��'2bh$���Y	���f��7g���'���M\V��������:ޜ<<�#T�\w���O�%��n�|7:]8�����N�t�=m�а���3�lTʑ�]���<����L&l��=Wv0� N���cypሔ����u��UyCƳX�ھvM�%���M���:E�'l�G��wnOnk����N�V<+�O�j\�5v�&E��T�O��͖!�-qF�u~�$x��eŞp�`iL�/}��ot��p�j?�=T~����c�%�����GYN�B� k���<��c�@ R�+�(
w��Y*��P�^���2mtMV��Ơ\���{���[��H1�3�_Z�nSU�g���7b�����`ߦȨ�%�N�{����DZ��߶�H�%�x����a�dԢ�.�e��S���3� 26�S�Ǐ�`֭o���f��~��\�����K��N(^�|����A�|Ǳ�[�ޔ�-�,f=W��+�u��s�{���?�c��P�}/]�w� FR�(�#�>i�~t��k�+��0������5kRzK�ٲ���0v���X��B(j8��/���T!b֦W�M�:Ҍ�8��61�ե;�jDq�)�*�nFZ��wrM�Vf�=� c	t ���^��jvΗH���h	eҖ.���V��b���?h2��-�z�v"���4N�_�~�e�Ù����H1��`��f���&ikP߈i��o�$��$����1-��K(�!��$��>؏k~I�	�_
�FO�^.�w~+�쵮4k�0�m$>W¥r�$�����Z�9�agU���/�Ӈp�L�2���Kc��'nP��A��Kn!��J���^��]ǝ�Q|�p��d��i��,l[�\�I�D�9��r��'c�1�	")�lyZBvv��%��V��P�>�ir^Omu�&yX�h�pA����wv���3��g�.�.^�q�H�[̙`�!�ݴ8:�.���D��B���%�"�")�����Sv�3#M�+��)�*�0��E��@*���VY�Đ>�>�I� 4�����n��rɋa6E���
'��$�x�7�Ɛh>ب
�~>R�Sk���r�Y��󅴔�֮��a�YS⦰m6��"��'��Wx�b^UUT�|%�@�HN�XQ�M0G��i��,��i�*肜��~�=G/�t�T�>���=-�{�3�����:��{ª�E��h��$/J�G�l?f�RP��?�4v��)OBd}��5c�R����wY;G�B1�,����n0�s��V�r`��*?���,ײ5�q�?-���u���n<�K�V��
3E�Ŵ�\�F�5O��}�WLһ�=~�i�t���_�i�[eǒ
�׃&ŶS�l հ�;����2�؅Z􇂮�ƀ�oo���j5Y��pQ�� T�ǸU�{8J�]4g���*��J�BcX]j���v����ف�XLK�cX�Ŀc���g�� ����[�%��A�_3o����"+6�7;ٞ �%TB ��R|����o��3��?��{W&P�c�C����Wm{�G�X3���i�r����ܰ3�)*b��˻�Um�}^)�D@3S�H��$i�����C)zF�7���T�Rϟ��ܽV>�r=C���5s"�����"�9�lHa��[�!u����u'2P�Z�m��1ƛV��.#�0p3[�飽מ�17���^L�=Ф�V��Xm�F�*�~VOKK��W�����-���ώ�T�׬n���e���L�~^аqTi���<#�9�tz�Iq�L�D�Np.\'g���	�?���ԥK%G�������3��$�3a�<K�L��%��6�v��O~9�hN�.�G__R�.�P�pH��Pl�d
�M��j�Z/��l�LkGV^��f0*�j[g��\tK+�Xr�0f�t�V�7��zR5��il�+1.�H�R����3)��ofeI�JF/�׼!��V��I�+gH�tJ��%�>�g��߸��h22t�!�Ҩ�������;��M�NE�vϒѶpA��t�=(5�mN>�V-�+���rC�7��HB�ļ��Û3<'&�YQ�s��2kc{�z��|���_�{`��ⶫ���kH�d�p�]���E�{��'_m�<�ң��.�c���oפZ;�;��*$<z��s��	��Y�\}v�V�c�d�Tp}�����h��bm�#��y.����_���	��+s�r�9��&�{����hm�8��\!�R%o�'	�v?�ޑ��:=K�jrA�_��vH�U�#ύD �PeqX����c�>�:#<�H��w�>��ԑ�p�]\#Q�S�|+x�8F�ٶ��$9���gF��N����	��_�eL��g�}I�^�ؽ
�ͮ��`�r������Q{} ��#����=��p��a5���s*�o8)k�TlW�U�c�=�ЈV�_Ѣ����k���T��%fE��Y��vA�u�4�X#���2��e"�Ԃ�Q���2D3�豅��'��P�MOƻ��}�<7\?��6Z@�h؊8�`���*�X��|�`�9>�E�ɖ���(��|��m:�CI"����p��oI�a��ﳰP_�);��,�Y���rZt��Ѭ�JXg>[B�I��x�K��'��Xx! -W���7���l�B�wc��]yF�g���& �/#�b!��.�|�d�������d��C_ڥ"�{����i�<��V��b�G�̙��HP�;��ed��o����Ζ��Qr����[�L�:�0�s�p�c���a����hL��4��^& ���g�[�����2*�YEdc��MOp8�y�`��t&qqM��9�1V�M����4����O�kg��s#��!�2�`H� ~.#fV[��j�0��uU1d^`��Q�A���ԅ�G�EU����߭Re
I)ddD�����g�����z�>�l[��R�C㻼�m�V�\d��Fм��>���_ڥgE,��@�4d���(�\��d���:e>k���&��V��v��@�a��5�P�a}k��u!\���4�N[� �P��f�}�#y.��8���"���w�%�� g:'��b���C�L5��RG��ه��SH�@W\���O���I�w./�ɠ-�յ�i��3+
��n�9kv�64���̭���d�O����^��۠���O�"/�r�����7��QD�m�{GF�!y���I��B�4N��H���7J�al����	a�� ��tz�@��x�8.fR�%Ea��45��oV������s}����6<��C���d� L5�y�+���D��0V;���I����{������[�R1`�/~S�k}��l����A[^��=n	Z\�����:����o͐5�Z���V���*� �QH�l���y��u�!ȵ:һ���n?0O��|�UZS��.����z!�f=x�G�h��֠>Wu����<P%�Ǆ��'�_�Sq����4�D�Ę�>,�]��6][gR�@}�+g4CG�(�UA�TL rEX�/&��H�\�>���L��G���J+�=J��?�7����l�k��Q��<�zgq��ߟr�f�8�6*,O��Ou�O�L�5~���I��Q����M�,����,�����xxU����?@���!]Fz T������b�qe��n�=G<�
g	��
�dM�������/�P�&��_�fJ���<�+,(;���/|xܹ�{���!��úUu&����kW���}���2��l��5�#���<?�1�zY�6��H4;�����_��.swL�(�\z��͑�!P�v�^n�b.u�!��������t����T�1����MN{ݨ�j�'������������.���xXY��e�D��d~��� ���9��<�ՠ�kM�¶�=������p���Vʵ:L��A�Y�sZ��lM�Q�|R{�����Y�=5���	�{��/�����^��E���un��hˌI�j�4�Tԑ�U���@~���/OZ��6b�R���8;�<ڮc"�Y�k�{�`w�k�y1G��*j6+��c�����.��`�9�!n:f6A� @���W+��:�Ld}E/�ǟ�ٔI��#~�y������vm�׹�)��Y���I�|w����vP�a��_�ۃ�m^��Wر1���(j�����[�;�<ݒ���pTJ:�8�`2l�S��0�Q�b=W�r�6k�-�_�	�{ҫWW
�Ë�m��^�Dh���Y��"�-`y��\���@��"��^�ճ<onK��L��gG+LUd8ٹX����A�H�,;�2$K�-���O3���&��iJ�%L@��Qс��n(ѾX-�b+�vÅ�U�EѩrQwK��'�?���0�phk�aK���Bp��Wd�
�I����
���т�g�{U�3�-+�������ʛ]ׁ�����4��O���EdĘ"�����EƠ��7Emc[~�W��}���2��;��i�����!*���(�b{���j�:k�s�0�X�uPc�1���-���uX��z����#���yE8Fa��2e:A��#�����f�#C�%gI�!6ߵ� XJ�����=�r�CT