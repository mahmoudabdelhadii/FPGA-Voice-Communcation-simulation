��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��,�y�}�ǰ�=4d�H���`I"��W�`r���T:tB�T4D�m�)�	1��I�t��
��8(�8t>s)ו�."[�漆���]�~�]��;�O(1#5�-� 偙O��QZ��~rL'�x[�i,mׇp���O�I43��4d�,�H�����SN��d���3���r��m���̨T�I;uj2Y� Er�*p�Q$Gm���p�V�`�2^���,hz�<p��l�Bxt�5��s��\yq���#�@W���f:m��T�	,*�񞭋����_��㧋l�	�\�:��uGd��PǷ��N�I��_����Tuv� ���us�(H�~�{2H�:Zor�Q	#%�3ˠ!��iS��95�,?�.���/�F�i{#���Tp5����Ҥ0{%���2vpn���X�����@l����3dc�ק�3	�Ed&3�ZN O���z��s�yxӡt��v*}ԫy nj#��lc��m戭k[��5)�A#�����8�!�]�Z�s�M���t��w�!��'ÒE�rv��Ϝ�c@<U��\tq+��&|�&X1)C�����r�A~��B�&�����s�:n{p��͠R�X⺂L^��R����c���f��J^?��ܣR�O 1�rV���:��T�4���AD����˩�F�w��)Dm�O�b,�a���1$��c��7t[i2>�ޔ0,S���󧇳Ϟ�ᒨ�-��}�!6��Jyv�醊�^_�(�H�(y^����o#����X��3-�k\8�M�T�"`R�DF6ȕ� �,5�;Ҭ C�k���1\������k�t־9�}���� ���QHF��"��t�9 ?��{E_�7��!����]���-�p^8�3 ��TLM��q�"��z�����`%F�zU��K�^�Y;FI�$�*,���!���w~D�A�]�#����u/��eס�yl:TJ�a�ȆJ?fgu��!0m�&��ݧ�g H
A�g�
��*����Թg
o���F��'�%Y2Q1@x6zm��S�u�ZP��i�mQ�o��=��,��n=?�M����j
o�k��MD�՝�]�X1�"<Q�}�ev�ߵ��Ŀ 	�ZI��R��c��Ro	�������.��k��k;7ˌ5�s�(nV�ZNe���O�}�y�f�����=�("8�Q�o��[_J����eUYb��[2�������g����-�������b*�̞�E��^*���������Y����y��A��Nk�j��q%���4a>A�fb=\���-)�����VU�ɜWE�'AH|�'��C��S#&[�+�k��RM�����rND&J'U��q�"C����e�#D	-���-�w)<J՘QY��E�~��͆.M�k��pt�%hg� �ྉ2�+��Z����]B�����X�K��+�JMDT�������<�L� �O"��y�N.
�Wn)bHl�%se �k̓��x�13p��~3`�	tZ����X/��ĵ8�,�6iԺ���v.�TE�7ҷO�{0g���DHDz%�2!2�[���i�C��Tx���r�R!��?Zg��,+ʂ6�'�36:�<�Z6�ٯA��O��m*T�Eu��D�gU&V�9+T**Ƽ�D�T�Kji��1A�2�RlkQa������*Vl}l�7GA�����Y��U5?u=5���o~/\�#X���op[^��3��դ�۰D�+� LmK?J�l��'�Ͳ�Pd��m�z��������	�=LX�6�2^�p����im�`_�=w�f�������Į�;X,�|�y�����t�t��߷O|;崰�^ �k�2ɳ�Z�E ��J��J��c���6�#c�FR�Z'ZvP,���E!S�~!�Q�1�	����1֓�̜�oZх,U���v ���Y�`[��IѰX��ӕU ��C̖֝�>k,G]���*�WU�|�J���II߉�#�'ݏYCN��.	�R�; ����W[�m��_I�ؽ����0%������7P�r�����2��7���E����`LP�p"MT�!?.�=}$N�ef\~Dү�$L;INf̋���UQ@N8ˢ�/.����G |!����2wr�
����k�3���s��s~a�G�_&�/9�դ�$�����zokI�h�"���]N$��%�%��y$�_�@��8�ǆ��}��&��Ș�邷�����Y��~]��ޜ�$#�I	�cqYхŮ�Qw=���Ǻ'����7iLX���ԓ��ξO���\���2x�}�I���J�dP�Eҥ �2��d�K4:�|l>i8��kj2o���(�f�| c��+ϐ�N��VO}��Z�9O�8��1�o.�L'd6^���7��&N#9�nuc
��N$	?ȹ9-���4� �D#�Cl��G�@;?�OrSl�Nj�d�$���f~e�9��xt����3�̖���	�\�J�0��AII[d�����JM�~s"J�y��F��ݘ�!5S�?8ק����9G��W+���ޢnL���Ĉ��ǋ���6d������d�W�>'L�iN\��f�$�tc	Q�:ⶎu�0ma�W]���fpt�3�K
=Wv�9��a2���%��y�ޟ����0������^�6�k�Z���&��>�Xϖ�l�=���e�R�Թ��dWj���g���^܄�<���~_l�*㧳����_���W����ެ�Ãh�r�J�nnn&7eIt
���,7�^?p�3�t�r8�J!H:�n}RF��&Ė%/8c�������*��qY�\9=��oN�Б1�a�;h5"����k����w�ý۹."���XR1z���z�5޳&�b�D"s�%u��S$��h�.aѬ�ڭ�?��fP���̪�/+���/�)-ևML�\���X�v�P7�g�����2�s}�tR���h�5jkA@�o���r��=P��4ٮ]�4��fH��k���"�P�R,���r�ky9�Ъ׿y�-zn�sӣol�(vC=�'����̆�tdLx&�A���u$�B̆yLR	1Q'*����x�|���e���<�ٸ� �_k+%��E�C�ގ���n׾��?P�i}ԁ ����>��ʦ���
����HP�)d�q�k�0@�3T+��֑١�B��΃�/v�:w���:|�\��m� ��n�&�j>����jSt�� ��@6f��ο{2�����.{9��4��/�j�ӷ�]
����PG�ce�v��� 3?/��0��?��k�妮s�EuG���?MHw�3�V���7Aha��p�߸b,�|(�S�n�4&���[����D�M~��2V� ���"��0y1�e>pd�=�a^`P��2�5��bC3����E I��<�79��z�`��z�" ����2�Ő<@t�/�1��t�Uc��㘇w���l��*�+�C~ol�d�(I�x���Y���C�@�f��� ;+]?�-
�EO���DknP���B\u��Oy����o��+�L�ɔع%)A�`�������1fƞ�v�X�5����,�g~�.-p�{�O%p�>ջ��IZ�_ܽ�	g�C�v���վL�<�q���9mێ��<����b0����~W�pD����{	E��0��t�m���;D�Ս�	*���}H'��vxP��cZ�95����N�p�z o���RS�qH��L(�-�9v��+@��^{k �Z!cE�a�1�l
�}#��hz)(rPAԟ���W�wR��~E ��R�S��'-y