LIBRARY ieee;
USE ieee.std_logic_1164.all;

PACKAGE bchp_auto_package IS

  constant poly_cores : positive := 1;
  constant poly_delay : positive := 61;
  constant poly_optimize : integer := 1;

END bchp_auto_package;


