��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���/�����Cc��<Nb��.�x{�>��0����=�����=8RLG�h+OLزV����ݗ�@��&�K��4cbXu�6@A��?��I�=��O�s=���
�S�i\��D���d3�q	��9/�I�w`W?ދ�S"K7��5�,l��C���
@E=D��!
����荾Z�V�h��c,Dt��&�����]4w9K_9O�=l�uE�w����[R�\�zÚ�-J�$����åCj�[�
����T=���K���h�����,������#�z~��?�G���B�~֨1)��k��yq�$/ju�YA9��SX�{@��mWt������w�F��r���������O)�mC�&�����$��^_��|�����=������A���_"�s���50��-�ݡ��kVE~�cu��'Ah%�����v2ݲK:|�g���7/��=Q�u�~��qC���
qSa�a�n�m(�]�h-�FK�]�Z<��K�b�s��'�����C$Yכֿ��h|�[@lXJ�*Qm?�аR��(�v�vlr�j)ڦ��0p�s�bv��jy�-����(��N�vהS��Y�n)!��\|9��;#�o:�#��9|TWL��L2=�'���$ƫ���19�?�:H�A���T秧���,rJ$�p}�a�ڡ�rn#9���~�1e�[e���!������{�T�7���O�z�������쉎�<o�j��D�7��lS�ƃ���F�V�:¦?�,�:4I~P�o6����2
�ԫ�#��G롔�qH���'> x������>I�nN1.�yφ�V�ǹW�)��	�3���k��c�Rw�buRA�8����\��L+p����rw3v�FF��8��Y��8p��s3jL&���9>��y�(r�I)ռ�I�|���Ն�[�.���ވ)��Uˡ�`�e�s�m��^-v��jEp�i�z�竺m�QC�����|��/ k�PpE��@��؊v���ڌT��\�b��nm��X�=x���y���	�����������
)���
��� ot�U�:�5�0���a֋���F��Ru��>���2��ٿ��V������sҨ�o��k�Fԕ��)JЎ���U����j���|	��|�����d��pE�P��>��w�P�������sZ2��"���<�U+4������r�T̶����M���ZX����ͣ��v�M(M�?57po��V����+�{XP�z��(դ�w�dQF`�D����L�y�*�=e{.�칹	)����C �m�SR3��������X���\`p�D��in�U��/�H�pu��O���M��̪TA� ��N�'�Q8�����m�\]2��P/�#tbFx�㲐�j6"���-���_e�HQ�qgf'�G2�F*��I�����\��D:�s!��+��9��e��~:�o��t�r��QV��R���abF��q���ˌ{p��I�!���,l�P�wL���@��鷹+)����c��<�X��)9$��8@��Q��2�b[���n ���qM�	Gje��\'r�a{]v��Gh��E��hݱ�l�O�ѿ�M�A�J%a�s<����J6d�dD<ځ����_�$�3��x��v�ϓ���|�r�l�w}K���H��U)�G����Jހ������]Ϻ��il̳K�-���$ZǯtB��t�ԑ8�Nx�V���4x���Z�uZ���3j�vZ�Sl�{�,�
���g8zb>H��b��YD����W4������JG)���(Y���ǔ� �;ߔG]a��_����:�Q�.�[��:f���ҫ:��vۜm�m�����X(Aƈ�Tm�����A��>�&�=�����B���m���Ҁ����C���HQ��;t���*_�����juO���P��-��95[D�e��@n2�,�>�2 �	Ux�(ѫ�W�+�]�E����;E�q���[8s�@<��sz�d;x���cZ,=��ִ�`�$�Ux��eMi:��H��"�,c�1�`�O���Z'vT�6�kX�?6�e�]/	����GK�Z��M��r��9�w-��g�9�RT��s�H
W�f'7Os�p����ږJSۄZ�nhDGzx��[_����ea !i��&9�.4�nǫW��jC���惿
ӌ��~�yK0!����@�[xg)�H���#�Q[W�R�c���r)�N�8->4�)YX�y����E���8;|�0	�	�7@+���#�/����5�u�q{�VۉKBVyzvr�FX��c�����!�Ӭ��>|�K�}�����&�����P�>���fŠw��t
�d):�*�_�8��F�C�7:t��V	$�z��f�z?���!ρu�}3�4���O���*�dVB3P��u8 q�D�9�"�RM+>N���B�yq���^��&�Q��݃�v�tU�7)o�!r�EW5Љ0�j�ԝVc]���v5�szi�,	~����`ÿb<1f�M��wl?��41ɇ5N�(�B�2�齋���`�S�H�m�E�?�;�G�J@I�� ��.��ڒ�����+�o?�'�W��<�
7t�����ۭy�3�ϖ7�X�n��:�)���R;�"����~�[�m�}f��NI����̹�w�z�GZ]�/�#a�yM�����x���V�I24\�|d��}G"� B��`,�T�p�C�ٷo�;�'D���i�����tAWc�����OM�f�h+�d�e�="�P��K��Z Y�|�QZ�y��8�H��Es�Q�!,_��k�t�p�{�N�j�'�v�&%�b�D���S=��avL��+C�'�K�x�xƖ7�j�Fr�^�M$ԙ�uNRW���9KN�E(,�w_�%���eO� ����<�����nik�d5��P��?fa�$k��!Z����z��^-?(��(˓�	&o�Q]���7B/k��P�"�Ԁ�<ZZ?�6�5D��2���ܫ�-'�$1<�7n\:wψz�j.���`��!��b*�@>��zhyAP�#:u�e���_������a��