��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��,�y�}�ǰ�=4d�H���`I"��W�`r���T:tB�T4D�m�)�	1��I�t��
��8(�8t>s)ו�."[�漆���]�~�]��;�O(1#5�-� 偙O��QZ��~rL'�x[�i,mׇp���O�I43��4d�,�H�����SN��d���3���r��m���̨T�I;uj2Y� Er�*p�Q$Gm���p�V�`�2^���,hz�<p��l�Bxt�5��s��\yq���#�@W���f:m��T�	,*�񞭋����_��㧋l�	�\�:��uGd��PǷ��N�I��_����Tuv� ���us�(H�~�{2H�:Zor�Q	#%�3ˠ!��iS��95�,?�.���/�F�i{#���Tp5����Ҥ0{%���2vpn���X�����@l����3dc�ק�3	�Ed&3�ZN O���z��s�yxӡt��v*}ԫy nj#��lc��m戭k[��5)�A#�����8�!�]�Z�s�M���t��w�!��'ÒE�rv��Ϝ�c@<U��\tq+��&|�&X1)C�����r�A~��B�&�����s�:n{p��͠R�X⺂L^��R����c���f��J^?��ܣR�O 1�rV���:��T�4���AD����˩�F�w��)Dm�O�b,�a���1$��c��7t[i2>�ޔ0,S���󧇳Ϟ�ᒨ�-��}�!6��Jyv�醊�^_�(�H�(y^����o#����X��3-�k\8�M�T�"`R�DF6ȕ� �,5�;Ҭ C�k���1\������k�t־9�}���� ���QHF��"��t�9 ?��{E_�7��!����](�S��0�q��w�9��=�i]�1�GʦȪc�W�XC�|�$��}q�6����zf(����լml�dz������*�eLD�*�,�m�]ہ6����D�Gw� �g��' A��)�m���b��ӎ���o�6ūvO��=�W�������}��	����z
��z�&�P�K#�^Qץ�_������&�)�ٺ���/��U���WX�wK³��4�d{B9/��&�	�d �Y ����6��-�X��o0O6K�-آ6�F�,H+B�*�5	��~��6�q�?T8F��Ýt��_Kf��b�Myz}���%�l���)�|��za�ӗ*���>Tk��EU�[��2�Lu�uU��=��L��Vn����$a�9�f~U=w��h�l��r�7eg�1���$��=?	)�Q��^��(�OɦǤѲu����u�r\QD��q�/�Z�/�uZ�!���KĻX���ɫ���X�����9d_p����g\��9hӍv�d&�����p���Nh��L����+3�z�w�����N�%���v�����7XrJ6=�(���9'_��_��!(�8�}�̎~ N�J �Ky@e^^���ށ^�$�`�Ē�p���R%��h���2�ۑe��=�'�� %����P�V`đ8���]��)|\�g!��N8��-*���I����BO�<Ft��9w`�#��ܷ������2�s�M/I��`�Ϋ߷�I�q�s���qs��N�ݙ���$N� ����f��&JF?[�c��3��� ���u% >�n`�%��QC�|Y g�&1=�WIx�ˏjY9 C��h�^Ǩk���_KTлi���Ăq��P�CBH��{�<���[�a[Ȥ/��O#F=sDI��2A��y���\K�c8���J�5�.����ÇE��i��V(Ed!$4�>yA�Y���*�ԏǽo3���M�;e:S�gʆ����/4s�oX��1)�h������D/P�\1�#��b���fA@?�B7Q�uH�r��@p���؁PR��$��\�L6zɽ�	$�b���Z�9P����S�P���7��Nj�A�r�s���A?������Ŕ��
�瀿F��Y������l�0�>��9�W4�E�T�U��t�})��$��S�	�g��������K�55�5������6h]�M�_�]�E$���cHC��=��SH|0E���p��ĭD��H������	w�xz�������t/k`z��in���"�,u"�q�Eu�����K�<�Gp��xA��f0���u9$��w�@���34�/�N��^�x��������&R�a����d�h_)l'���l�z�g`yP�<<�L]��?.��3�Ġ�Մݼ�#���_ ��;�cP�+c/8��M�:�O��!�l$ե��e��[Y` ��Ŗ��:x��H�yRB�T<W�M�q��#��$p���B�蕑b��/p�v7|N��~hz��6j�*��	8�)�Q�^Y�+�����P�d���xG�����b\����#���-�EBҺ��i�I���fIN�Ŋ%F
�8�R�ITF&����+��<�͌N��jṲ5b�x��K[�f�AO�eC��K����GMсA�f��^bL��0���7y��K1����&�|بI��T��0����}.�V}�?@�2�W%��lb���T6��a�8�2�v(H��H1^u}��`?@���D���YjE�f�!�]�t	:��L��0N��2x��D�ŜV���V5d��ň�N�{v0�TͶW7:*�	���ш^K�\ʾ�.����Z�Qs�=�^���\4Y�$��p���]���h��$:EL| ���fL��)�!nD�aT��s���J��!9���<��h�k
��Nol|��ȝaV�jӚ����U*�s^�ڿ6��&	c�9�ɽ�g�\����b�E��R����$�1���B��(���b��H�tt�%������X���Ô%���S�F��h�h�K|�Bp"��֋H��w�7����d�����z��y�M����1�H��=�i�4\���e��+��h9P��:��&����.L5UR�4Pt4\C��:Da8��G�J���^�x~9Vۿ�� #ۉ�Ә�!|�{.�~|�O�����.x���U��;;�M��(�v����D��+��0�b��$�Rf%����=oN6��:8�l������XЎ��q(�e1�5���pqAbK���ա�Ͻ}A �`*��'~j����F ��ե�C�u�.�$V�t2���t5����2@�QԲ��^yG ��5��K�q��m���G�{����e3�o"�?g�����;��c\�ĕD��k�M!�%_	�� ��T�i�f�wH�<��������%�R�s\j�8���#�������X]8|�J�[�����<�w��^Q�iL�]��|�H=v�µ���g�t@�T��xܲޚ�%�ܼ����[�j멝�3�f2S�KL��Է�K�0�U��)���"=�� F)z�9�hNͥ6�Z���dp��M?�csc3��])����K	�����͏D�!&&Kp5���h�ʾWĶByux�"�J'�u:~3�� ���W���c�eT���S�eÛ3L.&[��B����ȊƲ���RH�{�?�uf8��L@NPd� ��̭�c�P��Or�\9$��d�e ��
�<r���w$�J��c�!.h��<X�d�k��n`��H<�+>�X7:#����INvhe{>,8"?�PS���p�#�rOf�шB�ck�?�1�R"!��=�������%~PV2q�s7v�q�,�鬏~��/W�bZ���-J�M�-H�>�%쏊�%
GvW�I�9� w���]������m�=Z�T��=]\��/���/�M�yxyM+�.�J` �ߓ��Hq^lK#�lL����r�l�iFg�ß�gȿ��Q�{�qucҝݷ�ӊ٥x��b���*�uJ?�̏kHez�t�V9�����;x
#�i	�S��tf�j%z���L����V=� ��ˏI֎������<գ�>�2��r�	�|��5���� �㬶)�|I�<!���H�T5��Md��5�K���稰�h���]�	�(m#����g )'��
�[�-'���=&(�^�����62��U����Ux�G����lG��P�Vf^DfXeNyp���"co���TO-"��"��o}߃�B����wi?���,�7Q����o�ދW[��޶T_P�?�Ù��"^ƪ�1b��hm���\p�O���j���nWs�@/��*���	�������Z�+�鍌 ���!j�|�Ey�QD�y��PC��P��^K%;����<V�ޓ�^~�!��*J��h�%�� m	�w���x��r��8[{F�%6��3��[T87��6���-�u���*�#��n[�Byb�u�����L/�2�P/���0�ĺN:��I{����a�u��ZJ�.b��E�_Y��>�^^�v}�)G�3w3@�(��!�_�X����#�C�%�,���M�A��[	�p�tK��W�DH%�'h�L��_%K#U��c���v��@�5|\oIx�O@?��w$v
f���!�;*�!-;�JN>`O�0U�i�*�U�;ۚ�h�J�i!W��^�}��ˍl`�M��,R�.���ێ��b�9���N�0�~p̼�g|��%�u$n�h
�sW�{��~��N��T)� �6�c9o��}��N!�V2G��t��o�ę��m��OKLxqʜ�="���y�b��!X����;�<P���r�d��sKu(g�7E�(���]�9���*n����X�&Hmb��\�et������ַ_^��$���Wi4�#��S�P����En�z�B��:���N��p�k��2ﲓ�w����Y0=��e6�{��gGէ�F���Ɔ-�V�/�G�W�q�]�M�"��c�	xߊ�"#~FCJ��Cx����� "շ�x��
��|������ԁ�Ɔ��&���ؖ9�i�E�LQ�a~��&�f���(^�O�_Z����
~3��j4�KO��͔�'�^�E���V�U��;�q#�,r�nW���.Aאj�0����d�,q���y/��4�/ɱ�;,J#Χ(k���F���Rk'�T���� 0�;�?�3M t��:F��G��Ϲ�b2H^1'�/��bx��,1���*GW>A[t,Xג���d�p"\o�1$�&\�p�����jH 9�)�`��^=����{�|	��O�0�����9���,��Vw�s.��ay�z!�50�we�@����� mƲY�����^��x�B��� ��/+�Q���;X�b�m���0L8S%#�]7��k�q�����|�3 j��Mw%�U�ee��mG��,�e|�b�C���T���7x�w%F���2����C�`-�o�� [Ť���1C�O����:�l�鲠s拵�j�J�h�5H�L��������V�3-��.���]5�
�*���ڶ�����z�Vm��ʢ`����!�� ���q�ڡ[0���I��ˏQJ�=t�t�M�|���c�S�+�|�E��$xߊ�s5� =�N~�EN"헫�����w:���H��+>oi����aJ<�>1F�����Rɓ��D�I�r>��F}�;;d����[-S���T��n<�
'M�{cwߗ�/�5��>)=�\���Fحv:��2<�칚��ůq�ҌN��\�+�wBY�:�*c�I��z���m��6w��OU��a����>s��m�����k�!�u>C���N�)�(gc�z�����$�g��+�ٸ|���4�1��-&��s�1�:C��ř:��֓â��O*NCR��2G��E�VQ�^O��(� *Hi�X�(���T�~�ͭgm�9�R#�m�@A�S�&�d�4�n����xK�e/�Aو��:Ř��!�ﻔ�g��)�R�7����p��E�z�q�2����a���PJ�!+bu���0��u8H�S���Uo��{Ȗ�eQ�+��:G��J��j�o��[�fޗE��Eg]�n��l&4X@��RR��Aģ���#&Nm:���H���&�:]�+=����O�Zm0�ӻ�)�DW����=9n���&�-�B�8����,���rӂ��7[�]XK�,��)@��2Ml�K!t�|���|�eQ�� ��t�Gx��`�o�~�����t')�����U����@�-i�q:��t�| �ZoB��G�\RG)�as�n��'@5�=�b��1�Pi=뗉!�P���	n��v��yB�w�K��hx�U��HH��L�ew�m�P����[��x��_K��� �r�{-8���$��Xz�
�"%J��;�U�<�'��UI0X��T$�V���x0K� lF'�qEq�1��{].}�;ʠ�h��T���T�w&����ɱ���s���i7o����ͨ�6�ᦍ0�C0ADs�1�C�QP�������\T(���~�e<HF���C���'{�#hVHp+a!D#�k[+f�2P�w�w��K�q�G��B� 8�T����A�����N4�J�r��.l�m_~]6�ʭ&��?���x)B.s�﷉��Nڒ��y �UF�Lf���
�y!h��s񽴺���]������L�k:vl�rm��<�>�l��rB�i��!���{w���O��#�c�Du�x��&���H�;�ݭ���)�25 .9�J�C��a	�Pݔ�a�{���z�Y}�et�xV�~������ʬ������Ԣ�`����H3I�s���_o��Ê �A�@����d�3�R�#�a��JW�d�����2�F�l���Ď"@��ѕ�u���v�0�M ��[ؘ%�K�Hqs�������Eü���[�	�"���4�5L�R��,&�C�@���46���0�>�Y����N��u�TTq�@X'���ΜU���8��4�>5��G ��]��kLh%�g���ʎ5`�ӛ
1)J��I�M�/�?uO�ѝ�\�n�;���Z�����v�\9��p�ﬁ��Y�[�����[o*�_�eD�3r�^���_X9Ԍ��������q��@�q�c�����-�d��]�.���%c���O��A$�6m����#~��KH����w,�u?YȞ�8h����\JNU��n�,t#����Ǵ�OP(^z���̦�8{!hQ���)b�r,gT}cf�n�ә�ta�$��TT�2���	�O�	s������%鏁����3)4��WLnQ�՚;��������f�˻R�H��q���Tg�guJ���h����]�6�K|ԩs�%E	��^���w@�_�neW��JK"����W�h��t�S�P�����c����o�Q�l�/|Ʋ2�6;�>�-i1
�;���H]+���!6v�G+
9��u�2����_�c��қk���9Y��PA��\��QB2J���^e���o偻TKc��vg���y�ٛ�'J`̼R��7o`<���d�ٍ����SoEq�6m�9Eb��]��fH�����zğ�qFDU�5`xɧƐ��uR����y09�Pb$��^=����x�\P�X���zs-�}��Z�l�6�:�@!l��>�Wu�U<a������lR�-����Q��->���ֆ��!�Q� 6B�Y<^;sð�M���x@��`������j<h}������f�D��_��~���|�xė�Ai=�R��ꩪH��옎>?�Wݕ1 �&�D�"6%d���#�<@&�ň���I���wVr��F2�^��/�&��oM�9���N#���X�M�K��0V�������ډ�l��;���8��hZ9g̩�J荨�Q�CU�&���4�����L��nT$Eujg�h�6�eD ��H��C�GKc���z����@+��>}���6�O�P4
2��P�QDJ���C��2��A�q�KQe1�m��Z@ �|��ެ`x`����^�x���u�0xx�`���U��;����A�� 0��-�:KՖ��oG%T-6�v\S����w�DZ��`vR�� g������zr����@��gQ&m�)��{�E�����j��"p���"�)a��(���|C6~�N��B+Y��8�����M^�V_�5����w7dZȥA�2b���u��v��0�T��iS�0S؞��s����W�Ԓ����U og�+�ǔq�x��\z'�,��y B�!%�R"���]ld��J�N��.�	�޼.�B˦E��vȪ߁&�f?v� ��'�|o��g�����sX��rAì���A0Ol��k��u��H���;A�%tQ>�p��!>��5�������K,�6�ZZb?<���}��g��9Zub'�ǂ;$3����fg��=s�Aq��gM�"{���Q4���@��5I������ԱбtX:���X{yɐ%G[�E�	�~>� ��x�x=U��$V��tqy<F�e�kz�l��}���d9�HW�\i�ER���S�����Y�y/D�ȴ�E\ �Tl��8�u�f���	}��Q�jR�M�ܜ�U-�pأ��rS��g�.���\�o]�!l�t�;v5છ�˔b��|�����L8v�p,��`���ɍ0$o�Y��j`W<���!;p�뷟"�!��2��Hd�?G,\u�e5"R`3�iw���x\�Ds�_~����#p��0\��U፺�tn`��M�z\�=�?��JZ&nj�L1h�~���I����n�G��
ʵqJ vƔn�j�fĴ�9�z���?�:c�L���;��%��8S���G�f�������M#��`۞�Ȏ�cPq(���J�˙�1�o�$�*�X������n�$��f{��sş�X�����4w�Sx<����C�ߎ�9u:I�i��@�����m\�%N�B����5��ch�T4�HGG��kV�%�
.Iw]��ת�S��@E���[A�]w�3O���7G՟qJ� N^��BQ��q�T{�=܋�ϡFL���P�3�_�ì#mO��j��ڝ����­����K�����}��@IMt]~�`iz?A�i����QW.�ޥF0}����m���D�v �vw�KK06�0�t��5�Y0={�D�G߳����]��ƃ�3��Q�ԤD�# J�s�)�Z}K���ұ���'�*���r�#�G��j�۫v����3�:R�	�ҍ%9���n�4�)gA��
ʙ�ؤ@,w�\� d ��E�Q�t��o[S�ul���Pj??�F��<߻y�~l"�E9�y'�������C�7���I�mT7��%o*.��.���x���tf�i��k��Z��K��)��<���6��	�p�g�ߩ�'M5O�̌HK��hC��g�代���9�Ǩ���y�
���p�d�h3�9�>�����y�������w�0�ܚ����cn��'~�{v�d�����(��7� 4rS�� ��fɴ�y��]��V�P�� v+w�
8�b�7�D�Ujs�����&�-�d��S�[�_�o�w}�6�0|fKZ�U����I�(�<�e��`7�"��O'��9�՝�^�G���luI	9m�Ph��͑3U�~�@v��r�
|d����\�Vw��l]'W�2E��6�w��vM�肱(�sޛ�W�Ά�]�l��u|F��c�W�$�A����0M:��)]۪��8d��%�Y��
����0qٍ��;_]� �%gIx�
4X�q%�/���
��"ez�%�Q�����Ro�xZ���Z�g��D���2@�/Z�|Vj�8;�3X���ur�9�['8s\����Vķ��a�;Ҷ}���'W���G�ƧO�<����]�֍p_��߃?��gx���z�����o/a�b�[��d%؁�I��akFGb��?ޕ����f �Ż����Lզ_�r. _�O�B1�˟)�;���2m�1��_J]8�C��*@�R��ai7�B9Jp�o�����X�r�R�鮍�c^qށ������p�j��xNH���G�m��>��mR�O�\g��W��g�.�H�2���q�S�K�8�\�3;g��q���U�kl�9������ ������I���!r�S� 	��WD��c�zL+Q]�S��ID�@ULD<d� xs�Q^kL9�J�/Ɖ�M�:~. �s�����w�t���tLg���~麿�y�)���l�!~c�X;�S�t"����(U�����4�u���s�$��n�͚no�ޮ�3@�T�f����:�e�sP>�鳞z����y[\�i�o	nj�B��c_jZ�LK��襆���r�c ��>K1"�|)�b4�<��a��I�uG���~��R��t|oI:��~�g���s���!9(O���NHA�TF.f%(��F�G�Q�A�L��p��	���Xd�1|p�OA�RVe�$+���>�(��Ay���b:�|?�h{`,?��F��@b-��\˭R8B�M�7=�rk�l�*��?�v�3sRs�cν����wO�~z��[DKE��R��׻��O{e�d|%Y\�������&�䪃�En��I�a9�b:n+�u���u2���w[�E�.1�NZe� G?�Î?�\��
-2(�����y"�0��p�8�%��~�Z�x<��r����h{զ�L.>ꋤ��u�fsQש�����Z����oE��S�6r�p���-�����N�{�'�;�=[=q�QǪ;_���'��[�W����_n&E"��0�]��/ql3�����?$�X ��I�������S��J�̝#v���>	jf�J��O<��D6J|:�yV�+ ҟ�~v	&�9�A����=�L����ϒ�6�����ٝ4�.�̇���+�}~�ϖN��<�xe|ڡ�9w��=<b��mQH��@�YgW?	}j6�<U-E�~	5���g����?�U��/� >���A��-׭��+6nN�\�w}�B%�P���G�Z7�j��# �5zET�y�"�5��u���K�5��W��dt�_[��ɽ�iO�)U&�ſ�ZW�UH��u�d��l�t�8c�sNո��5�e���g����gĉ��:3&:������h�A@�;��5�a��>1|���e������|���uS�/����صTu�N��������[�o-�fyLՀK)r���u9��N��'C]7�cѨ^�e0�)T�'o����U1�-N��U��������~	8�w�)��nT�i���M@�"RR]�;�;hY�4��%�����N!��zݢ�5fu��$���іvh;C���o�~�F�;�EVG�p�RM���3���v�*�/�� @+��Fx7�UEߠ�1`)�.8t{��7	�4l�K�.:
Rt���;����=�@��Eu
��Z�z�GvH�\��oDLU��YW������ٹ  Ϧ�д���YY,Mu�c�S��O�[2[���*���L��u�//Odv�i�Ҥ�\9dh#���s���O�{;�K�!y]��ԕ'���� ;V�·�����W�hI����r<?��ij����,1���x�G �ަ����<��)'���Z��w8Ў�Zi�6�χ�	β(�l��>�DCՊ(�d.cA��0z���k�r���Ȁ+L��F>��P����X�+��&}#L�v��]Ij�k� �����j�����q?:��'�`'��0 �w	�jx�1O	�x�g'�l ]�����r�X����/�� � E)a��[r�N�7��z;*1� �(ρ9h�o����Ύ9^����~&�j
=����	!xV�M�ա_�¨������b�������%99�P����nǏ� 7�AL�T*Hc_��V1G�~$�;�(�-ДjE\@�
�1���sI5��`$�����Py�B��L�!"׋L�IW&�E�>��״��`[��ʈ4��-��)��P��g;��w}$1��uPgzh�<a���R�u	/	�
�f+�Yݤ��f�,���sT��h~$�.o���\X"�ۯqݝxr!M��X���-�?s��9,�W����2��&T���G����.�Q���˿H�l�]�F���]�ͬ厙pmʧ��U:eX�o,J���CɳR���.ߕ�-q��|b��i$�G�vI�4M���'�c��3��V��,%��4�*�Hl�	���q�f�L�􁬈Q{�2�O&��A�^�;6���H�FHb�
Y];����/\'Z������ ��%�XO��x�n�)��d���;��)#�,�2E���㖙���Y�̟a��H�_�g����������Y\O����v6���� s�&|���T��Fι�T�/��i�3�O��V�HC=�2�1_�U��G��hOS><.YxZ��c�{�?���ҕM�7�Y��������\a6n��{�@���:�J�M�#f�NUn� ��'����A��!��Őa'���n��},yx�/� ?�rG�hj��`��}"�K��O4}��|��Hv��[ґ���X����ْW���*��}���;ߋ�������x<�����(z��3,�A��O+iґI�ȋY1��������F9LD.�@HPb�s��d+ba �Fd������'�q��S�C���E3UrfxP��'M(Lel�ઐ���>��m&�B�x- Y�w6��J��4�:��cV�0��ڣ��1]Y�x�ײ���Kr7sa�Y)xϮ�M�O�b�=�̇>��
r���b�+$��������hhv#��FK���׶E��,|⃯�����>�	�|�yϑ\���O�NJ�.��!y6�%�Z�@<�����.�u�^�!���a������L��+�.da�R�S�Ft�/
�}#�ѷ>���6��1�?Fs��\�Q�x�n��	�� ~(e�Z�ڇ(SmRd��MĈ��/w��g�P�d�b2MTBx.��3�����1�����|p-vL��%� ��P�rv������p�'q�w�r�i�]r\$a���O�<H�f��ٮ��2+�6�|I4����v��vJ���	�r.\��r��s���}t��B�$��_�z\V`٭�t�*�&�Y.���/�yM�
8��R���n`�S�*��m��Q#Ať���E��'�y����$�/�He�J�O�S�."
��]�q�aؚ�W}�p	���f.��B<A)z��lG����k�Ǯ��I�o�Sь�Dˠ9�n�_��ۃ�O� $����ǚ3E��=�?�`g!�v}�t�k�Ё�Z�.)�?����U��������?J>������S�M�5������,V���h�r�z��4�8���kT���3F��`�c,uT�>\�^>����hҋ�	��&g8�i�J�4�_!��j��[Tk�V4�Jj?��p��.؇�J�4SC����}y3\�!������-���d�l��\Ho /��#$<gR����������]���dUj���bv9�2P��m�`�	j���9� �?|���^�~YZ���R�'��w�B�.�W����l"�y���}�8�h�W�/1�}Cp,�*�:U�1-�� |G[Hs��Y�A����n��~�5f2'������am������"0:��L�Q����|��P���0Ds����+:P/؄�".3������bzPwZ��JUӲ���-O/F���(7Q������ oV��N��p���Nu�,=r���~q���W:裉F3�X�z�y��7�m>���KPQ�X����3:�;��{Bޛ�N��}��QC*{���ad-��~��8=x���-�S��?n�O��g�0u�}�����-f	�N�3�u��0F Wi��d��Y��#΍j3_g[V i@#���M�[��T{F����ҕ��f��+�``���� (0�X�:Ï�}\z��Y���{4�:`5[z_X�r�ꥠ0����LTā����5?2� ⃗�M$���r�)�S��5�W�f+�;����
�V�F���,'/5EUt��ɚ��(�j�ԫN�/�r�>p����.J������#��{	��@��"'ѩx���C�vk��1�['�
�	�٥�W���A`����ߢU���Yp�]����:��N;4�(�%^��P�x{��c���W�hT&�:X>c���hN&)��Eٵtu<���)��Z2?�r9h�/	<���������:b-�����a�L�n��|����Lf3xx�^K��𽇷=���&��H��Q���E���$��Í���qC�'�׾��t�~���ɍ�[�� �	��?�>0/!a�B����$W�6�-�ʲR�̫�s�qm�v�V	h!%��a>��]C� �(�B<r��ʹCn������U���F��M���NEP�^��饬���x�3�O�7ϵ�5��8(m���ԛ����t��5��6��9��SR�2�3�ݍ]��t������j�^6��z��A�r^V�S�]�+�2�ڰ3a�t�� ����w�E�C�-�zP4��E���
�k���E8��}R�&�4���Y�/۳�XRj����(טU�R��Z��3۷�fZ֛�tՌ]I�O}�0��@���Z4��܌d�!wJF��P���ʍ��V��H�I�	l�Х����r�3�h��9_�d�Br_����ًǙ���u\����3�o�����dv"�YI/�nY����fȽs������ku��'7]g�#4_bz���x�����(�r跧$2%�3_�D�_E1�����Y��6�3J�����s��jV����}� �,X�g��C?O��m%��/��ve�l����s/�7@�Q�3
�ͦ!�m���Kʫe�3�+^��l~6V �O,b�i>3S�Ǳ{�("���:	d6����:w�G��F��i�8qϵ׃~��EdЊ�� ����d�ěe�^i��u���?=�R$�A����rp��fi�
w�=�0Y��0S��rI5�/3�x�� [ꄔdF���qo^u�I��=��ƪ�"n���@Y[٢w&��_<3�H��Q�h�Ks�h������C��P]���"ٗŶ禞�R$C�ʔ��a�����fVX�ʄo�b���2��T*U���ܚ}�A`4��o��M_�q�
0X9��oi�_S�39�ij���LUl���u�:�J�͑�p��z��-qslLa^$��	vߊЫ#�L�e^���[�-�G!ϑ��(�R��K��=W:���F#��{eEmv��Z��ɐ�ʛ�w�pO���I��/�+�<�,#b~���a����#��E����2b�x����=�(Z�Q���Is��#�n�����I
� �
	�������*���כ\uR�d8����)��E�(�mv���X��%�!<��b�_t@��gv�O��POZr�P3��H^����+�sNE#S}bM�� %��>�1�0����W��9
2��_�]����W��ar����ű�I�II�_��q�Vs��"A��غҐ6+m�T0����&���5��A5��F'��\�����kw�i�b����e�NX*?�j=�_X��X��>���^T���"v�?W�Q��J���~�#��?,��e���KB�������̾��Q�	�\ձ[�<M#9j\Mu&☹jC��5;��I��(���������(6�#�`����)?۾ � 3���U�a�v0����P������P��*	уf;%��!�K�.eͼ��`����{>qc	�.Z�?��h��~Ҍ��n*�����7�Y��
�"�E�˅��R���c�N�ο?��gR���2���5�7*�,,˸����#m%7Fuͦ�~�`b�B�"��U�$gӇ�G�W!��<��?`��f'.¤�K�Es��X1��te�+�QJ�@H�a�&�t��
���Z�D@Z;`��V/"^��v��?�d1�Zȶ��9�,%���#�V� �f#Ci3�������Ɍ�r�j����%�0��Y�9Q����|v�����/|"�@�'=紐P0´�b��.��P0�^xud�,Y��omru$ɦ+�\������¢�O� HW ]g���<�&�Pρ�j%
��f~,�(�g%"y煠�-znW1 F�9��Y��#�آ�L�f����bר/�z���:�}�'�s(�L�~�f5��,�W�(�L

�B���;�>�3�+�	t{�쉂 f��"z���o�� ���_������~O�(fӇ��S�P�S�+�Rn��8�S���\�����]2n���7y�^���=ѳ%X�{�E|x��5�+��D��`Lx��H��{�l�u�.s�=�� ���15���|��N/�mB��v�*_�|�Fy��ĕ8vy�aN�喵?���J��x��Ԭ�a�*X$P�wl󊜌���AAe.9�b޾;�A�"Ag4Q-��A��%?�pN�7i$R]h��~P^�H�>�A����]�d��gֵ��Q�\C����؃]��h�TA�𽄾�X�C
p?��ϫ��ߕsL�
\WK����a�{L�G��}t�굪ۣU�~���XXm:�����ɤۡ�Ia
,ſ�L���@�r8��ტ�Pt�|A^ɨd;F~r���G�1���r���j�����B94H�O��@k�5�n�����c� 0H���&D�f��=�D�ӏ����e�[z����W�f�5'�8����[݉�^s��x�iՄ	��;"��}�k:2�p�j��Dv��æx���ށ�B��	��i��|�>Z�[l+ �HO�4����'Ä���v����j�
��0ߜ�BHf"J��w#��}�'(�֛��PS]7=�s���6�z���n��v*&E�aD�gX^.��'�ݤPgR�r�3��1A�����FP�pS���#���W1kp�4�+:��h�
?�T�6�l�����)�	v� �x4��x��@���2r{PP2?��J:�'�b�w��Jju	7vk²�d�I�v�k���M�@VS��j�� Ww1k���l�e���A3�y~��������������r�އ���'r=��_Ƣ��΍}b}Rj��g��~���V��b����k����9�{$Ż��T��o��XL!h<�1w<Z:i�����5
�kp�����[�8����ç�K���B�yH����;0/K�'�luEZ�V4��W�����ۦn�Ј���60nu������nc؏K��}��*�S���`Yv
x_�l�IF��}��>�k�L.��������=;����{�L\H8�[��[���z���6�SmUqsO��9����-=of��S�_�@���ye#�l��5��B��b�NLI��ɄY�G�ɝp�].�Bjhd�� =Ľ�J:��g$�"(l�n���kL�A^[�Ӱ�TDr1<U��N'���G1��6�	t��\r��K��U#WM���29����k;:��$�li?N_>�SE&���S��LO>�����6p� C��1�pu�3�V;�ۡq��)�_�G ��"�W"+n�p�=�O�P�uDx-^�հWuCG�����Œ����5�.���q��j���3�*7k��;l�tr7#H�B��Eh�;�<V�� *����^x0�'����5҈�\3��z�1�'�����T���y���u7���h�7�75J]����]/m� Ȧ\�R�m��%*]�|���ߞ���	����j���MH�%��E�e�P�Θ����}z�eX&:*�����@���u�9@x,&��Wt�Y�?v[�-01b��;	�RÚ�Ho"�E�[��B���%��>_/��~�ߪ����郯^;���y*��I$��>�l����E?zb��&Xr3J��8�1�̏$��~�ye2�����J�0¬u0�|k3��<F��S1�W) 3�YG�	R&jfI!Q��h�4��4�x� �@	�ɢ�N��2���'�B�yҿj]�R��)�\��R@(��Q�D	慧�/K	���x|�cQ�Qe�+9
�6u|� �����W� X6,�i2�r>��:V��Ou7Z��ɢ >���9G3;nZ���v��u���o,-uWQを1-���:@L�I����e�|�P�)`���;8L�k��9[�[v?��Z���O$�.����?����CY^ij�e����e�kh�蔏�hp�����M�hk��q~��;ϑ�f��=�S�7��5rk�V�y����		����ڬ��X��&�0*fd��E�`y��,S��"�(�S�t*��؂�W�_�;�f�cW��nTڏ���f�n�.<(���r��0��W�g){v���\�jh�挜}�>�����F��rk,�d����ꊙ�N����W��H�`�,h�j�Ԥy�iB����:X�`��vAE,O��E��H�e�޺��/�v� &��6u!TkpX_R �K5h�wŮ@4 �-�N�Q6f�Ū=}�M��{0eW5p:�@������?-mܺ`��8��	�T^&��D┡�>�T|��p̤����kK�¡L�Y?-�P�{y�wa�󄻽Pn۳O܍sy����_V�H��rZP�yύe�c���|9�Ꮰ*b����;>����B��Twks��\��Ļ��7��٪�~����/6&��u�1�..7"�^	ͤ6����'���0�<��r �ߛ�0�[\%#�f��T����>�h��o�(N-������w� 2�_jߋ�ը%�{�=˪��<c0�Z�۬�/��C{T�a��$����
Q�M܁#��Ĩ}ˬB�2i%�3��=6B�����7;9��Jg0�`��"S*�{�Զ>G��~T���*о��R�|�h��5R-c��X�I�9r�O\��ꊕw%�ve�&�P_2�xJH��7j���ůc	������f27�I����.70�.�͔qT��R*E��eC�6�[�D��q���L��6�9��������JĂ���o�ap��?��FV�^�A�x��i2(ĭ��=�`�B,��e䖹$7aBd(�X�����s�+݁�EM%e��2fԛf��/�o���8߫V���|���q.�L�	��������Ng]ج��UtE̷�Z#�n��b(#�X	o��1J#H[��e���
�2 ��ct�f����Y������L[�rf����T�֝h���m4��`�PZ�!��_;�F��&���2<0:�㶱����P@z�2�2��W�m�h��&�9�s�eds�ks�Kw�Y�7��e�8���J,�S�D �R���x���N�[$ƕ��0�U�~[V��Xs�f+��z*f�"{{���S�9�uM��K��Rf�)�ݨ�df�7s
?��C��n�T!�m�Ÿ��Uڒ�t����E��
�cI��t4.��4&���Z���݄���L�P�fR_#��:FW���4,(��>}�#�m�9�|WTH�����,F�O�0I���_�T�-����q��&wI`'����l�޶4�4��
O����Y��g�~�5�e�yߌB�x��v�1�i� �tx-g��h���&GZI�+p��2��QcUK�a���x$��<Q%dk�<aF'�Bs<b�`�E���6V�!�W���5~�f�m