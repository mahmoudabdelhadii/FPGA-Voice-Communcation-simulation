��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��,�y�}�ǰ�=4d�H���`I"��W�`r���T:tB�T4D�m�)�	1��I�t��
��8(�8t>s)ו�."[�漆���]�~�]��;�O(1#5�-� 偙O��QZ��~rL'�x[�i,mׇp���O�I43��4d�,�H�����SN��d���3���r��m���̨T�I;uj2Y� Er�*p�Q$Gm���p�V�`�2^���,hz�<p��l�Bxt�5��s��\yq���#�@W���f:m��T�	,*�񞭋����_��㧋l�	�\�:��uGd��PǷ��N�I��_����Tuv� ���us�(H�~�{2H�:Zor�Q	#%�3ˠ!��iS��95�,?�.���/�F�i{#���Tp5����Ҥ0{%���2vpn���X�����@l����3dc�ק�3	�Ed&3�ZN O���z��s�yxӡt��v*}ԫy nj#��lc��m戭k[��5)�A#�����8�!�]�Z�s�M���t��w�!��'ÒE�rv��Ϝ�c@<U��\tq+��&|�&X1)C�����r�A~��B�&�����s�:n{p��͠R�X⺂L^��R����c���f��J^?��ܣR�O 1�rV���:��T�4���AD����˩�F�w��)Dm�O�b,�a���1$��c��7t[i2>�ޔ0,S���󧇳Ϟ�ᒨ�-��}�!6��Jyv�醊�^_�(�H�(y^����o#����X��3-�k\8�M�T�"`R�DF6ȕ� �,5�;Ҭ C�k���1\������k�t־9�}���� ���QHF��"��t�9 ?��{E_�7��!����](�S��0�q��w�9��=�i]�1�GʦȪc�W�XC�|�$��}q�6����zf(����լml�dz������*�eLD�*�,�m�]ہ6����D�Gw� �g��' A��)�m���b��ӎ���o�6ūvO��=�W�������}��	����z
��z�&�P�K#�^Qץ�_������&�)�ٺ�u#uD�	' �/|�qf�M&P)�tL�x�?�u�����ҽ�����*c"q/�\��YDl2n֢�vtX��Q������ǰ�6K�gVL��ο��Q�������-�˚e��"gb�_� L01�D��ثU�8-��Nw�@�$[�>V,���6�����=����{>G6��v�����φ+Y��	�d�A��b<�)��Gp���k�(�vWu����!5�^; :F)H�	�>��_���c��'�dǃ~d����.��2I�$ �m�~���/�A.��Foꨊd�[j8,���3ʔ�V����4��VT�����V���ujz�P�����!�M�}j�eN����Dt��2����J��i���!f�[�k����H��*$�����*� ��Ɍɓ����>ao߫�Z�Jؔ,1����0M�b ����cEf/��R��}�&`Ԉb���rp1@�Q����h1Ci���]����A|�n�D�I1�@�t	�eɮu ���-�`Xd�i�u�\?�f�{c��^�߳a���ZPs,tg%��2p �~�~���<��T���u�Fq ת�-�N"&�0�s.M�q�P>��՝�P%gN��w�
��fD���k�cM��W��Ժ!���8�� چ���T7�"i�Υ�S�h?k:���c��JiTg<�2ʬ�TL��MX��Wk��/��N�`lQGr%c�fk�؉2��!�P���V}��'c�����|ۖ���:?�AM5�3u��6M�]�&�$��i��ڕ��Ɩ*������M=Z�,�s;4wxϴyґ1ӱ������D_8f:Z�~=�c�]oe�-�h��,-�L�>z�O�T��2��GS:��8.��S��	I���]^R�����8�~�F[F�w��/g!ݹ@G2��	1w%۠:�(�A�[�5wY�{b����8��F���~�\��d%e5R�.�y���q�f
LG*4�Y�b����Jd�=}�lI5Ŧ{��<�$��ȤCOdt�Դ�eu�"�� D�]�!����z�CH^�!h%�z-vR�B_����4��}����	�Y
Y+��E�AQ��
t�'��j�w:gT���a�&t�ך�K�r�]���"?���O�,N�Z� |iJ���ur
;O����,.���K�+S��yDU�����)y;�.�Kp~'�g��ን��rV3I8����Z���,	�J=��Ş�nVs��/�0����ˬ
j�IO��|��QS^J�>L3�b�L��(.���f���vj~x?Q��nBP�