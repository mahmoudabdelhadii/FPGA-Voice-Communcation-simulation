// (C) 2001-2016 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
qRjY2BJlqY0RDCP01R5CBVkrKxUaEKEfrpJrizr97Kd+dnJxt1q5eCngr3SRVuohnkGbjeWYn1Gd
n0paoyvHpizU9PPazItt9LV0ulJiGpGyyVXyx3FR/8CpJfKsYEfcj8A23CvxuqA87Ey2/1g+q/0F
pnxfX+P3lRCIUgVo15UfM/g/9SAVN0Kj1vNogtOiPbmdoC4LmXWe3pKLwXUSxS328Nesz7J7tCyz
VWXRF/6P5VmvNTUFLIrLkqdUy6FnVcUKVKyGqiAsYPLYOlSWi1b3T8q9tGhRaf/lSOpKEP3bGU/z
Txlu3wxSe55XJc0Ys0CgvlBUd1GOU5hsm2oEBQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 7872)
iAJkfYpp1rTT0xLzcxzDvBM+NlQchvcKQw6iz5F5kQLr2D54MvOfNk6ubmGjrY3owa3XS7RLhN2Q
VC9ESahXPEH4CwhuFHNd2U6NXOGHAjjvHctniOMUh7pvkL20xO3GHIJA+v4rE8q1UwSNYxPudZck
FJ31q60s1Crx96NweqWtWYSyKzH/YfUTN0VIBOIOCtqVdTbX5C3we2MCr9nRkcLY+giTuu2d6OUy
UzB9vJuskoBwJN9lG42l3XWP+azPmN9xope8B9sDO2tXp5uW9eC/+1MF5jL9TmUAhEskiEjSRpkn
mmkAnZ49kIoAsEolxy0+sXmU/k5a7Mj9SuHQ1Gl2nnr5DNVC02fSquDB7iH24177T8THoE/3YLQM
9gwbphzZSxsIJFYzCoZ+31xSstNptn6v/jJxn+I64M3mzdPZuK5gsAQ3FDBFcgAPjSM+fOTxZ+XM
rJse6oQot8hEZFJPX1FlVAN1styNGvcjDYm58lOD73v6Y8QDqxUQvPpZLy8NkyX8W0Ebv+tansuz
eDohQ86zTlM/ca7lnfLkeM5OS2paAwIFX00547bOK6kfwgBilSVi3FDeECkIMqemz8IRMz+dYSkF
p5dvoSNew782m4H0lkAdv1J0iAj3YqnC/5tN+b++DBMB5jhKaRg0FZVHhIhRi589b5smT+EDeygS
4kmtoAuv9FTiLQJJLhKRuwQOn3AIAhNw4QwEk7wJYQqBrxZkTTmtugwRrrmM3SCDKdr7M03TWgLf
pVrsD3AT4fQkYYdH20l+PrIZTtaWly8WnxURMQYQ/OpjLB4dokTb3d8QA3ZuVzoW/Kdhu24fPcon
MrU7aW6OVRJV8HTY4aficl+w+uwG+kiNFDChpFca3T8tBC6kH37RxSjJ5LGwR06qYxj2pMDINqoZ
Ay2XkqIUPPGmkbxFZ73vSDIx9ztTLSCLNevcdi39uj/M856BA5SejoUAjeKzhQiv9RiTI+7ubE6D
x0QbE/mYE5DO0tvWBf+EXlMG6dBAa85Q9xS3txKsJQzZLnujzsUKAl+AXmntT8esoUwwdXvy0wEz
WTrOZF3xRdxqVz0tK8zO6mB3ormM5qwuvj8H44IQTFRebUOsDuqaZZphZIr/S3eaAuxA8cXQjTfr
L8duBzQpYMAF7ns11UkuRKINoP6AxMUP/YrKAYIair2k4+KW1KZGhMNbCz5lc1EYly0zPw6LLnX8
dWi0kjF9gMdAgmUFndOMahwZZ9Xb/025nVgQyBnow5WeCfCOD2u3VXs2FEYvPxTXVI5u/GbaNLU0
9FqUnfRGEZ7RDvoNMKAF7IYi4o0YSHDscspBbV86Q9Ut1IAmwvBFnzv9ec19lFq+7xeCvVcn0r/+
jnxQjDzjaQ5KFY4/qMfqvdsGbY1UWYzFAwJo8TpLI4NZ+O3HvKAJcA3g5tYVE37nt9q343XuHGcp
7S/JhM1gXg/XhqAFziBMTpaOpLaO+hrK+jGxVaokwX+SkrhYsly1u43NGeEWdyBDlrwI8g/iOoww
aHLvS4XRmFnZ2ygMl9MKZtw0TuxwscYnXCX6tqh44IbfIg3myMy6lePN+9T+RI6qQpQDK7mhVYGD
seTShdSDRricFyoGOf2PkL+qraGjs2zm46DXPfFjNmffWW1CbZj7OKY4+LWetbJbhfePXWVQhpw8
MoPjZ4Q+Vbv8LVW5670mNkivzqCI6JWweAWfIgpKsGeibr3xgZtBKpnllae7at4Hhm9aEHQjz2jq
i0glC04P/JCRwuPyhp+BYI78p7Zln3tY8ItqHEOCz6zVIcaiA4wbFZOeKCV0dshEN0Y7VwE+V/be
8OUEFf7n6GweWkOiaU81VKRohljwl2YP6aKUIN5zf9HNVxu21cHzNVZWa/xhbT+Y/T5lgkL4ZcOj
vtyCrhNikq07P0Y7NDQjGn7DRlgL4i78zMuKyTYq1nIh05b7Yvkk2rwdy78aO8aXitz1O9PGW1pz
TowyjJk/56CKRffN/aeC9+kEd/Jme+bERFF+Lq7LHPQ9qwA9QkhUUOKnJZIeN4EENqMRqx80ZKrt
1/LFHKv/KNWHtyqQUccjkxhp4I3x0lZ1F3lAQHSQvUA2Kb+Qf/HIn0IfuXSGFT6/ui1DVcizN9bD
RJRAUIENRC8nz+QUtlzGv9qE0JPARNwwpDVfrBuuel+SuiqHnkzLnIht4Hb7crDbKgmelHqCXS25
PBXdRDa7GecrOUIlnm+7JZVPfA7hMnCFTYA9jGWn13UMbcMD8WkRwPrLq4Mxg3p7eTBF+JB2SnRU
ngeA6PV29rCKQODdVnRIK6+p4KIDqOrf1BBgy+lkBNyIX5rpQUOPjWV8B2cnV8WxfVfQ0pBIEGzu
hhWJJA3j3ceFrHF9gE++5bB1gi2pcQysGjyDPT8fxCZHUFbm2GCr4R1P2Qs6UsM4/O7S5hFERXiP
idJlCWJkQ45swMNmSl3uOObj1XpwiMKNEOtFa+dfqLR8k/ZWFx2HXxQd5jEy1YzBqXB826dOZIpe
28pLiYEXg0ogkETTyFUqtsAI4u8f6mGYYDOqlISyXIfMrTZon3PpxUioP7bDqr3XpDW9EN7EV6aq
MffEK/KHbi/cNCMbgkSabTprHljlqF3jxA+Bs+eAo6xnuvG0OwgEbskzMMP0I6VXrSYebBm6teJQ
aKAqaACUSYpY3dfsMFO3uBvJFOYLKyoupeeggmp9Xxoih9u28ohH/rU2liuwjJXoLkZyyzTLF5RP
B0rbZWJxdLe21pXiQrn1fdadgz7EFZRN8RgHakgunDu37+UNIrOAIN4C6vkdU16bCgB6LCbI4uke
QVTfCAvlJIBZ9itTCdiubO4NHHCM0avKxx/exBEoAuNZvBBIwXT73jJQhsfswZiUcr8To3WGtPO8
sVLRvfgwVj5eMWrjiSMfsPQrZPpqplkEoPTzgDsTpOr0d1Nr8rCOzytfJT7+iuVztuUhzGYZzywz
G6++W5m8kmbWtnaMLqQG/gvVzYHxyulUlRILEz1QjRaIcMnM5AQLkFerU3n0wqwM/LQVpVa1WhmA
wIyTPWGlYbXxUu3OyiDC6nxdXlhaks5tCcJfJNAzBAHdLKAw+iPwK+738O7Ici1Ti7CZfKmKc3OE
prse51xO4Q43ri606OuEtn7MgBjZ/wG2jh/hvZ6X0hLkupWauOFh3CNJ0hgOQl4OuRS5q882dBVp
UjRkRbJhq8YeSMHBliBYd82FVQatf9pJi0iTv1d/RpwL2Xi1XsKKYhBPsXtRRKSLTIIl6fVYEzaZ
vAW4aIC3IGezSeHXZgGWN2Ldhq05ylAwUohp8LvC1q7c6TqyI1yEueR1E4KP6hcHMjlrLDbu2oN4
bLZRGPXM7Dswb0DASxGnYyLsV8S7u2SkilHvXL/Cj01jgs9pztUKyEcDdymSQE2+x5XAF0/hv88B
mURiaxP1PMpFUUdZPiDSf8Gdy6el7wn6KgrBkA/Ea0SDOE89mS9Fi7BmtyRKg7Hl+7p5Os2WxNCd
ruml6Q/qD8VbLjVIRRxxbzIODRpl4HJ7xsjt08DDOjg/A2g43zDukFGCe45WcBeksGwn1qplgRJE
bZKlPZOSMkmshIr5pYaX0hjsq+PwXWk5iAOJmptceoozYPUDPh+eowPF+nWFQob0O1pEYV7uL1CP
j7EYziiXyzcpCOYbtb+YZJeBhG6H5TbxTEkuZ0w4FGPvF9XyE3HboEytvyF1ElutMuQM4yg5CS1I
S2dyEr8KfocMnL7VXKciTUsY5MaCqlc1IToCEDPJNmc88hugbETbIQ3YTeOXIe8W7q6I8MV+s7R6
TqoPWrbb+ttAEMnowVDZwfoWqnGw12RsARIZ71esShZZ5lkplJoGhWiZ4mzb/dFJihdfhTvwW5Yd
Sc11fF/qRFiPeoeL4swSVBvOT3TVLCet2vtn2qbZNfxZ8Llfr7T1Dsr1+KSou8HzG8J0INsoIoR+
P5sIEIehGpbER//xx7pts1NSRqmOobLBKMJCS7Ui6YPVnSBE24qwA2Hp0H2Aomlw9EjC8WW1L/iW
Ys5TqMs1DTTzfGauKz+pzTmKM8D25sS15+ifYNFTs0/uUQALkqVxC5rJEph0Ry+IjrL9Rk92pzSU
4kIVfEweWtZUKt4j2AvSIQeLR6H42XCCmUwCXyLZx+Ri9IRhOgCM9ILdnWVflFdm7r4StsYcGCwr
Ub2aiBCENnRAP+HuVuzrU+0hq+wbSptpOdLN8VrYYL/tBhoBOGlZ5AaUK65O7WIiFduZVgxP5Cks
dc95IbnXYFKA/7pkEKQPoImoxfV8/JVZo/sHRWdCCJZ9SIjNilZhjTmB1tJ6RpOLc49Zv9cp3Y0d
hq3/6TSpAP7yQyV2jk1SSHyHZu98i415Hc5AQ7pXdcE4zUwvQGVO/297R+2YaMPTYuqOo//v0nP8
mrysNUBS0BwGGrY4BGWLHjnDFTQXP/aschafkPZXU/+ocKBXAyLJ0sYVcNUlu1+rW1GVZDF8UmO5
5a6TLBqLjRXb28t7xdxvh7gWSKkmRAO2xpnxFkld5oEaGrxsN7nHnbDH/11NK0px2v95Vo0Nw57u
Oa9rhPuu4wOc8UX/SU0JqnQcdGetC46wkuO0s3Ic3MHNVqDQqcUlABHQ6HIUk6fECiAYXlsD/PDq
hda78V2WNhMRKjat7V5WSlBXak4uV41A+pj4nhW4y2SWNSa1tg0hrxru/212g1wQns413lCBYAXm
496ZgeA4a7brC7L0uBz5XOz7kstw3PbBPb66yHqN62ekbvpbsfm1zvZLKQmDrTpY/gBacgdEBESo
XtazSdXhb8BTp7Wlvul1BKvXCR73ilFngZmyNA9oSf9dgt0rLUfXkaKKl8mlygGYesEX/7NxOfQ3
UqtbtcGrZjFq/SKXRDIJesalxIkPTO+HtPvVWHLDH9foWzJk/Jc0zi3c42eowAQugnpMb8HleB2k
UZ82twE+i/OlTG2gpyXyMxR3QBZUnLEhuWDE+KcD1aet+30rT7y7I4AkjL4VW8Mk6p75HEX+1qDY
JmwziyJ/j3uzaQ6Vt1RFlF8Bx0FjYMPbCM6/JHCz/ej7ahmZg2Xio4ptSbuYqLkfyCLDDg6xLIed
J0/M67hs2IhUsZMeclO8UEcLEgmo5Hxulc6j7dfUsmdGCILP7/s50kdaQDJZH1Oic8cL65SMZWzk
xWvw4Gmh/cOuS1fsMzCjexCCzYCfhCB4Zb+XCULh90jBsdw8zpAzF3A2UdptYoaMerqYvFNpoQUV
jGJLKFZCFGW84l8Fn20KGRdQUoC9D+TXBlkmkgtHOMzb15J4zHEwhM4TQ6qAwr6z8d9Gtyl1Z8wY
SujLaxirZ1RUs1ZgF4GvwjSulIlv1WVxsLN7Ty7QZ5jVZOGtnbR59k0isgP50uSYkqu8IoXPHcQU
taGzP6bgFlf/WRmkZqmRyxQM8WSm6euqNPYqXSYCC4NAAluGPgU7UQR9Vk6fHn8rUuIlVlB166Jz
L3vB+LOjqU3CGruYrtfOQrz1Bvu9B52idy+tZaLbpCOcEmnzOfUFo1apJ83u97QOnrqWMMNyEnSt
NbJ/JZ0dFJ9jlYuwgCG2qP6HEFeI5TSJnBHwQYAkbt48qANN3nCzq1pyERTQcfNKe9cDqpmK3ZeX
qBBF0LcIPRr5ClvYDwQLsNoAfS0xfnSvvT0Xbzv/BV6O6lJRFIKBalH2C+CZUGdlkE5P3OvKbzwQ
HhJyPxcJz0AMMGq2CGnV1rF8ovfSNGGTDaMyciWW+iJh/NTfdPVwNojZFR9vqWo5yraBrYT0lVBY
sf59bxo0YmH4s+jdWdrLPbbhFBQuAc44mnG1DT7aOrq6aTAQFrYN2v0aKAxUcC6ni+HkxGjmPLiF
lCVaMm8mbmvTNbVd9mp4EjYNBfN0FI0tygTRk1OzIN3TZqe8DNKoeoY8fbcdNFYF5pKGjlc4+OWN
6tAlwagdmy/vQR9+j75Q1FRUbVuCiqcTCYXS24bXnzuzotsx5DMBVKnJJpixhnPuMFrtTrl+vFq1
V3lXPanKr3CjT0/r8yoFi0R6+uUwHh80YQyeHNO9m5rzYDORRk/gKqNGmtW6tQQv17k/SbfxmnM1
q8bPwFnGxW2dCENF8UxSHFgfRdIlpRkcwwQcXvZMPm6nXRz/nPKirmH8u2qhMOCe9NaxnXHGcbih
26S3IcyVWZzkflBwolxFgaN5lplOmguXjJ4nHzpS5rLbomtTCg85K1MUdDCaPmz9nEqROxat3IlM
uJGIdiY/7Hn+CDD6Vnla03j2TUp40p6N0yB+OKVdFYC7GH9buTmDNfYUsqooSAypCMk//dyaI3Va
h4xY2/88Se4wc2aVO1FiCBth4XqQv702DzfnkQ4lC4SzHdjMLptQyhsCCVzumD4p9xHbh5Qya+jM
httV4fUvYKM0lRQV6DphQxeC0FskCwhfMicfOnuPXlqObpyWHyHoHvgtO/Y/12e0fIvjnbVpz8S9
aHx/xLP7FChDLeEQhCjQFbomd4n8qEDpileW0pMOgY5RM16shfiAByC4T4al2x5nMchkMEkY0Jei
5lsZR4966TsJcXZuwzA5acUbLnDMWYOzlyBLbFwr7JHtCeOQFkEOfM33re+YvEt2m+65mbmyD/4r
UGOkmL/FAHkJSoXWtLBkZbG+EJLl5Wo8EkCMbjNA6osoxmC6S18QbYTGODHuTg/xiL42zPGq8q1U
1GKpOG3aa34SeUwzrYc1ygKWUjaglvghrf+pNCyLFIXRccTecnBQWiahq0pn/2nyrK/kYf0q6mSJ
JHWvgfic87bSGmYuWvefp1cmAm/9rTVrog7HdTBbl2tgdBHM7vRwGwPTbtMdI6Pn0nc8IbKyZqV8
jbCZoAvVtNPkAfLBt6Z+s+EV3fqTnVbhWqIP/X4izsbU5LcFoeyEuJDimgW8RYvxVI5IdVWXZ9RH
EhgbBv8EGLD2aZBS1O2uBG1FuQl1s/mXESYTzCIw+MI8uSszqQFF2NwRfGfF0/J/v36NmbWHdjae
yUS5raRACNsmhJQck5DTP7e2sJuJPDUICgx5gOlntSOlGJvJtIwU95h3cbwguWD9Ph8ERsp8Fzm9
pW2ifkcTRNlPhfDVTPP7ee2cueECnD1iOPtxUaLHi7MG/0wMfwarum862UI7g223rnd4W+ZyzS5K
bWrgpDoOQr3PE36Jm7B322jxErLFfg3hZgTSLDVxr6K8CHT5VS+y1XK9Jzymf7iWX1N36eGftZAq
q2h/4z7vdWfKmBcTq6WgPT4GyDzbi1lsdeXcd8Zpw1IX5ZIl0GjjXWsjIPthFs9wT8Fs/1eyn4fE
zAu8YqO+vS8Jdqn4tDmVoPkuAg5CwQDt3GuLL9stP83u9Ifm0T5MSD06nNfBDV6r8CE1k3cUnkTU
P+1JdJzsxA2uUFKSaVeSqHur40C2kzCX9T7FPQ4b5DDVLBPgpdaajFZGHSEKf/Q43hpgNqfhYBOh
G4vF1C0QGbMhg5vry6zju+ifKXCdol8IcwUa3L5SHnncMgyaKfWGdwvEpDKvW/QReSGvBz6QFz5z
p46/T/ZLBtPhhnCK2I9IhDvY+peNtdJFq8KIRBHSEFB0q8i1VHZmuWLX8/tVGA6AHISgknN1bx1s
+fzdxZpPGNkAELldZ94yrVBJ9QHqrgZ0yESd1zjVn3R47tQBv/vGG8tcWnnnXbSvo84+PfAl13Qp
qou0Tg2mLjdTQTEBl29T3gaCJUKe60OLubN8P5f+SIwPdCUdMD8xRiOGsDJ4gKr8bI1jz8FH5fZJ
g/a1rOc9ILIT5Oj5weqS1JtrRAx2s7/+9KiCUOZVWHbDmeUyt90kVKlit6PtHW1x9V+Rgm8Akj/w
ETdKw5B03dyLstotQvDRsSUSR7J1mTtVP6wZAjRwjq8VvkbM7sXYgWr6tibUX8h3JeOioeosxJHv
GKx+M19ITXRCyArihFL5h2OI77r/K/3pV7WUHceXZfRxZX6rMVflx2E85yspC2FqpiliEBCnXBIN
JHOd+lEb7TajKtGGY+cjFT1lKlL7geZA9Q81DyUfeaKXRjNHHWUEVWydlUB5cqCbsCk5xG52xL8p
krGidwQ8O0xji0p2RuZgaXbCrZG/dqahHFx9OxYuMn6ZpinZe1M46tXsMGZALqfTCGkM9Obhl1Le
Bdc9lMkDyeWTaAzgQui4bC4nthEBjZ27hrDraaAfwchGSXhjJNqR1T644Ex5FNWpUn71BuDa2HiQ
fk1ejRrUbrxkloJtAfaBTI6N+qY8jdApu7r4LakbAyQt5YWtvEuTvjuA21fdgwTEHyTYYgWKx5Ok
k6HCzxAUSrxJZFiFzo8EaCodxCjzx8hcRCSCZ34AHOlbww6AITYrlXt/bEx+XgIQpDnHOo50sYIM
Aby3RmaOO5amIlGeHP07muZ25r2xoN33B7/ESF7152/g0gSRWx3fLsp9E+YbQkOKij8cBFvTjs4M
aqtFlWzKZCGa/w3uix0fr5x4HmulXzA4E89Ee/rl/9HTW686U8dumAeSsUk8WLt/++o/gO6zteSn
uUt1XZ1mdSdKm/zLVslx0CmoHC5rJ/hYfNXq6m7Mtc9/vweXHSd7f8HGzOGzas9VP6ADZZFOaMNp
ReEbSgXucODEnSCucq0nxc1r5qoB6rh5A++WhTXOr0kinAbi7EBkGfiO8+W5AZrFDzle1ufw8w1/
8oON0VAdOBRxZ48ALNFSca76Qoqf+ceKxwg2dB6f1oYQu7f2F8K1kseIqew44hWaghBNuwU5H/YN
q9an1LUNLdeDCwHaVJmV5tET52geYuQtMb4WLYyFC5GgicWTyGfl56Y71isXNQOMSYVKsH6WAT65
ib9zqE4sGWP/M4s07KboJwwWDS5bsq9M1pjKy15D6prTUrfXtnw4zIrgNLbdesix6p2xL7oqjRYt
+2Nggi6ll4+HAfQV9is8wH3PiEfBOmpG+nio/xCqSIq5J0qBIDfM1T8S6AcPUEDkSyQzeyq16FHF
4txPw6lw/kJS2rKsiRNmoDgGBgL4L6/YZL8R5yzhl/Cn3RVs2LHLraq73z92QU5pXs/o9XnIisyP
CoeJAtayEyuvK+M5CwPOpemAP3wyCEmiERa4EZXUmUpeZ8Ad4Yl+4Rb4DkLU51rePjVXNLfyzqJU
0ahfFxp+vM7DNrbLgR66uxfw9OXS/LmrRcyrg0SfZt8FIcP5mvuXFeg+g2aixRzGQqlxTS5/PCFV
PQLlNP3dYGYMlAIFoEGldF7KpPJ7lOUe4Qx5tjflvtDWyax3p7GlWKc4A5BXAN9EvYgydtENRlbl
baKl4UYGBBCNdsM8sggUs/rXaH1gv9jB1Rx7My4hnm3Yrq4AolUzNZvMq39fS/RpWrSFVkckOByC
7dTkUGst0Ep4tFNGIg1tCvt/2wzwfnyK2C8OC5HnTrP2xn87H2c6mHlBKQFbrOipuWwO7fC0BBd/
CStTdwxgGsGZCKH+/VynlSbSGptzuN63Qs1N/Fp12mdHfJsBvOKH6d3cHMFsgHCYOKCrby2O2zxp
680omNjDRsq3ctExlS3V2kaqfM1CadUI2GUsOpNshbCGexyD5ii6WfR85zbV06lIMa5bMlJGrAKH
ocLu0vE3bbps/LD3FrN9l5Su6lN6pPt1XUDZv+BJotg9AXUOnL2GEp6wbcMyIlhFv6Wroz0zxSBx
4+neRzFVdagfYx9qFpZ545zY7JoGpXo0eUqrmgemFZ5yf5hNgdOlYPpkLFXzDxVatjJ2kvMPNDu2
cSyMIPFXqWGWlb9WSyiaKNqk284J2r1IvQ+76HXrRyq6qW9FksqFYq2CUQSbUne/ZddSrQkaQeFH
X8PgZZGiigaCJZiXdsxAqqG8Sa/lmZ9olbboatPyJl3UogXd8YhjVZ9vdSGbqtM1vIq7CZfgsK4z
PQaICpEBMKJty9MbcIjpeA7Zt4kSQEEW9sJ57EbYsSPNsIm1JOtybWvPDTNxIc4rbPc9GyL1sr3A
DMJxc2HszF9mw95u+JPjlr+JY1IgPuRcdHgVidVO5xFFtJ5p08M7JU8DLaY6uaHQoKQhCBqOa9Zf
Kp030QwbVj9cLxSHy6S7M7n4yR4xSnmo7mPbat5AGxjT2uV8Dn60CbkNq7OwzY7fK0sN4H4JM5Hx
sCmMsPrLaE37yrhlQhNghWn0tF76jKDeIO6zeMxx1SLZ3zRTkk3m22AI/D7x+J4/WKNw25e8t9E/
mOWoWjYxbS7zzaeYxPLC7nAi+Z0eXrQq4JqGdVOu/9F2ak9Dq8/3ORU4DWdmWarVrfYP61T0M95a
oiRyQIpfNID4vgmsYVVxfiih7PLqd+dY8TkdLZCsaFAuq4UMyf9YdA+GfM83W7uUKeMfpGIeO9ai
VPVDC0HG1G/U9OA9AWUSQeaP4ReiDnQ5sfPfdSmSjFWIfL0P5VId/OaB1IaWheNSdUanUkW2+P9r
rZwNkAEC6d7szUPKlHfQkwCqwZ/ep1SKKlhRjBVceAs4qRCqC3ANOWFltwjA5ZWXMJmRbZrmA7iM
GiiARQmx
`pragma protect end_protected
