-- (C) 2001-2016 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
kaim45R8i1K4bYFCNUW0y+XqwzuiJEpSVV5jDz3EEHb5m1ZO7PvIcFu6DpbHYGl5dF39FncqPC7V
9s948gWesC9FSz5KIiBUE4SUB2fkqia9b1vkOSK4cLNGjnZZBF+ch4p41zCvT1wQvnHimedeYxU9
/a7wQ5zpLBXX8gD73OIctW9EsjpgN+hpDeI/ank0Syg8uqov7PXL+fB5LMOR8RPkUytyFZ6tfuot
ELwv3WHXULMf533YvsKRt3hMkmn7BTi7vsKDigw1PAnM0CJaeAAIhqiaHUJ4i6P5YJ2JAdkRVBhk
4cqTrpDHvVFFIpucwS5k6jwNzvDR+ASNcNv+Sg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 5856)
`protect data_block
+09ojmwqKQmw+DHARwIyock1zkgr74s1qK37jtapM1K8WWR+If+72gXvNNRhHQfsILAhAIdRkLKd
DRbuSXK2OyH1cWk1KKuOhvMe2nlzIF3m2xomEkBZdlBiWVfYjnfs6jz4/TOJ9qtnQZaIJoCTgNGH
3PFl8q4FZIc6Nm6N9zZpCra58wvIgfmSEKwtTxophB9Y/vIyuaYerOXu1vrr44Q30YMtikqtBxPA
eoRT1FHgdA8H6zx5nneYWQxzlNWOPDMsNeIOuLNfe8dCSskiSPeLgDW6sZL2DJrgU7i7eaOMMbbW
sPJ2zaS9v7qvlZFdQGx9vIMWsoUiGdpQbvhU0wyeb644iglUA6FwnaRUoHPhQRbTtwmycjhjz6Be
yWtW1R6IB1TG9EoE/Xh4Xiu7S8tQPBUOwaVIhbiFX68fYDPvYUlqE4EPU+JpPYL16yFyJH8l4689
E+EewdUXOxvEg5QmFxVK09JiWwFkFt6B5GsaI7Bq7l7tSTz/Bpfy2MkxGVcmZ34ukiBIcS3lXYrw
/HejXXM2YnzBA9vxjx5cu2Fbd9+WNDxUHaxUfVPiUhDNb1AIw4UyG1dw8yPtdjUh873laatKKX+G
XOF78jXRloko8Gks9XyJfr7jG93ol+tVMKKyzbAua3Ke4xixV5cNFoLcSBJKOTZv31vOuad5Q1Ef
5Keqghr3CLEVM7jTnOdnMOA8DsKt1h1p1k1PFCVuQ0tiiKh5+tGygJk04Hvqu468xAlAHvtET2aC
eiuuvKlOgPlw+55irhKLFczGSKVr45Uvsm2PuSgk1GxFOswAZM5D+OqJdB9O0GZ4pZrhxc1XYfWR
8qb3gW9U+o0YKApwKSFUCwoTOObbZHYaYH6kVnvax2eLAYVNHpAvodS/nF9AgijHacxf/JeEPx/z
jFyQpo9QAnQLpkKFhE5EnwhQr26B1Yy+qOTfjE352zSLg5AJvDT7NB8Bopz9olrJkJVBuaY1CQlV
DBQJWU5hUT3jPeIEXwCzbUHp5GzWuKew/dlTyvJcTr+xMM1QyIQcNmSMarsxkIQNbzcqmuI9oHXy
pRCbTWBgoGGH+nzj5mNSUYHuNLXYy2X8rTPpRWbMjYUh+N1OzHGUhVuSF08o0a3eFy3Nq4z+P3em
jZE6iE8KD4WkZopaPK0Z3SiV2GTlZmFYXV0DfMo+Ud/4xEL2dkgK9y3a4Q4Rpmz3T19kGOQdPeX8
A4HdaTv3geFUPOwh1sAApkkGmjqlqqSf7zQMJxqePULOtoyoGqOS2CH9CwrZabXTrC1tSEYwMDPp
KNbkXqW8iQOcrOTonf9YyG28jaf1aSRFHBVh6P6SXuH3Fh4jpEkYafDM5GsxZbopvsFMrWbRW1SG
O0maIYjHQs+5POoLaapB5Hhb45MP3IbCfoGo1hz151GMnaFAl0bdThciRbknnCTzt2B4U+TpOkWz
ZIuCkJRzf2XMDssJ0R+cVAx714kTnAv3aLvgSXldDNb/BEL9ckc5nBABq9tDIFoj1vZQNUGpBtwR
rCzpAaKAabIhcKW5CampXAkn0KlYNR7vBHAHcVDkqh/o7MUIc1zzR/T1kq/FS+UUjD8A042ENjS0
QzQUKTL1MQnBwQvon+zsW5ER8iq2pVlDjf4N0vYqwmes+6Xa5jpBv6C+osHQYfmYcpFyG3hN34b6
QTTf+h97WW8AP+YLAiRIVVxXMaYk9lKJsalcQsH36hfODuFwMeG0nkhipG3sgFCnBfSjFl5NjtGn
z9ir4XWqLgw8hilFCoglmHxhmYHH1xGLdP7K/kdJuRuoUWMN2Ri4pMQP4KrUUTwvMnk0ry3diDnA
COeGpYmjmf4uCvOWTujlKzb6mJg/RfZPQZpsPt2vqRQDdj1cQW1cWuvJghQ2y1vU4TDzUlOOT389
R6B+DTD1w5JizMH9RaMhRxAKiXHbx31feqkOkj78IZ3jYuQsQIDHxv/OgPb0M+3IRijwITxh+gD8
k5zGwd4iX6GT0dG9NswVGBIQfsdsQvSg0ML07l4MgkS4TmGgDXXnhWZ8AcwezMld7NG/EH3Ve8Wj
dFPvSZBu1VP0AcBt1SRGY24+0Sg2dggC2lycPjtX+tQRSQFoDHZr/6mpelQwTAG68CvLsaBjjz0W
Ntc2yZBVNS41qhRrmMy4ivoKKqcXhZeSuCLJ5N5lZ+EJbf3idiqOjY+TCe/eBVVdCoIlDBjNRTYU
jRpbKBaTXuVXUvad5FQMS1IZDh9tEVYhqKf64WT97ESWlABI/427QXX+I2lOv3nEgvGjxRG7E1PJ
P3+BX3S1QFkP5rY3iBsAA6bHOrh1anDKQdP1eV60t2Te1Y987p1oxWv7YEhFrE/M95/GBouNmXGj
Kbw0fdeeags2yeP66bj78Il5ZfBxhgxllu59T08Mz+EZhfiEtq96SKzIMpwWEuQipSnJb1RLWZrT
+odmNCc1QxezGcjSotY15A0uZbURfrlumdmXtPbfKAM2szaw+k/ACKkkRSuZcmZ75HRK+ybVbbO8
1BrRQ1+M+TM0hMPCi5k9Poelg4gW/Wi5nNQldcdUQSUpvj2vvrIOjyWITz7ljDS/mEgvCI/BycLE
IgCGVDGFbEpklDYKzC0PpMXHbHjIAjt14d/iJLcNYBtkssNZrT9XazqdpwN1t+4tng2K8tkGCCZz
iBznd/+7quUsXzSAmIUtgPqxQi+Mn58OlgWSpm2qdbvQZo8liy2nvyFbYbMtbl4C1wTYLM/kQGBR
s+Msyb/6czmYsTihpSI1FwnFI5C5FMHov6+I0lX2OfBLqSj6q4bmaBkWl31u7DO0KUGBT9E12sKZ
4xSIhrD2K5uoF8ZJfsjkA/ZxvKJ4oPBOUJW4PzcGFkJ72VMzfP03f/d+MuCyadcG4RZunmdRo/LY
32NETqqqpoHtgXGrFaO89ir+5kISytncVPEXmj6BTWfA3f8X8ti+PLwqhg81/IU5+JiKwwY0tEIg
0dk0lgZRSCMdcT9e6gEaIC7Vsjbd2lpxYLLpFXP+fZViqrYFKIcMNw8xMofCZ8SjOf+/DSLIAJnI
yi1Wh7bTxGiswE3ReumfX0hFOEQSCaJoqCbOfiVx5zIoYB6vURzNtT4loqXMrAFbcoRkqjjM0c8F
KSz/uaq5t2aoFVSPTZFLBEJAUIzOiXDtRrHTT62YlY5g6o7PVmU21tKx5wZOevY/7qi9woVCLh05
ivH8tCaEuFR2uy9ykpnsWQmqadeqe4Gdt6KoqLo8Lg5haZJBvJdEl7gtzXBjtp4ykkIRz/HwBp1X
i0m87FNeulqW75GT40aa9CNdNnxYTNZV6nkG4xKSLzDxX0HxxWgDp32Of0qlwNMlI/nkBY1+PBmB
mCuSjGGe98dNzT4UDtN3W18HAWfxrYj28KerjsBVSMDjbk9jBuxuujeTXTNoyPBoOk0ZmekmSkRV
EHY4xGo8l9C1olRggPGA6F3zLweCZmzaQY/RdfkHPSxzqtVwIAbfOzBKxpkIFYiPTRgytGmqApG3
JxXmWBQaY/YgQ6t6CBAvvLWfQzCfNf7Zlx8jAxgLYy+nWp3xH2KPTo3MP9AlFMYk9IZREV42Bb7Z
A7+yhuGVAkOLpp75ANdp/BTr1aZFPLVUmKneF+mJLRAuAbefEs1Ve3Ew6UONFCs/d0tQkdVtk4w2
etlt506LnRm97ga1IfBqd4ksWNOgR9OTLJh2Xk4X9opdSsRMua4wNmo2Lz0uf6Ky3zcnCd4IlBxO
Qzr8NFdgcx8dgajXhU7UTym783u2l2jEpSaO3Iq38c39cH6g1DhmPTm2ShaC4yOn/zSYx+whhpKN
fALzmxzIUBHDt4oWOmbsnzNvCK7ai4RBhQpWhQ9YK5AhCEljHUfazwJqTDZJGnnHoykwssX6Tdx4
X+OPKcDmeG1tTj+BDvzM0e0fA5OK6cHPbEBxJ3VEO9fQIoIayYP6eYEBN2u7j6f0g4jfFRA4Abvs
/ra04Llw7qo1t0fHva28jdTqnCq3Iqp3WVueUI/mx4M0dwlC6AzUiMNQgyml/lobsVY6V8wP30ce
hyUktQBGTcE5aCSHMbsWEYK9tbyw7p0bYvCwZAb6962FfzkY9gmC75XJMR10UkQKyWDBETAMUZPZ
kTO1TGrGnqZAflW6do4sHmG1mvAC2X7fOxmRwFtGeIA1S0hVuYbo8txNfj++GtkaKRBvg6EF75yp
7pCwYzGvuH6333c1w60q6c11sQfr49+GjGupKtwO44X8eUpCIuQrK1JWWKz3Q1cP8HZTdvPS53q2
GD2R+zWKfNzFLhtrfIrWjo2u6uO9lUO/bvuruCRWONyxLXTASOl6JElvR/0EfvT/5kebTyx4EaBx
GkVRRf51a9kHfKkhJp2bXReZgMLKfhk9/sQk1G7Il8tOYpOFRzwEw0D9vdqWmGf+a2tQjjAgTC11
qh/y8nqDwXVI3ArAKPlH8ix/DVdMd1YmfwWzbmMGV5RSy9DWwUNTrJ0RFFdF1qD7peHhLmxeU2tl
rbet29sXArst9ojqljxw+1mAKBFudQ4epgrejpz02ycPGHLSKVjOvBm2rYuDFajPAveDCmHa6vW0
lb+AhPrBbBdzr7tC7WKgNUnBJpzpQuvydO8/RkH/HBDb67FqbeKgcFV2RaPU7xR/BnMy0ts5WjuC
/95W0FZltOuIVjdfos1Z0wbEu3VwVaC3cDu+LgKCFXIh/pKxz/5Z9zbJlnhY4ULDDARjNab15V4K
9nWlPvwQj723I6YUt4TvOtcXNGRuflM7FHSEO4Sdg9Na5YEo1xVqdajh7PHdHIRPlqxjHHQPKnzF
xvf4u7MvXA+3po2RR57fmC/QlRa9c+QMvik2rPbzQ1+n//aPp9qu3F1u1r/u8XvS40GiSVmj0lS7
5FWgw7SuufQNYVkQHlRUrrbP2IH/PnxpowRyQZgwVidFHhu/LeFlLXlA29kPK/2GkEBAmBb7nozx
Z9JtHFbi41a72awYKdDc3FVyCHa/MdHa3M/3JxtD2Sv818JmQn7IswFL67Wh8rzv4Pycthps0SKX
1nCQzJ0eL3jKRKT+XFTKkM+zZCruY6bbnFnx654RpnXBciZZ3J3zr3Ep4JntjOsmwjREPi2Ccaip
YvF9hl2velqltUsE2Xp16odq6HW1D/gVRlpaAUjeaQRv9xPcuOVvouO6qzHneSVvW1G4ei/j3jGm
ZMPt3K6TFZ81qNDu+H5zJWkkga5syluwi96iLVQhhasL319h8uuomaZBmHPoiiEDcvDjCRPiLtVg
CRBNQmH8Knp25Ua2bOg3qsKC4DZBe3+C1uQ+iz0c0M+Aqm3yp+CMQ2m0Tvye0rQKH4ZakwyZOJrX
PqJjKuq9JgWp0GhdPCz5Jl+c9vn48m9T7h7XFbfE6HBOLBOlhqpXjoOOC9KRD1//m31KOKDarBmp
zoGYZRCc11PfYSEPwQuWZOqKY+T1xkIr47mTdK8sBnu2EDzoCQeYio0JGid6ER4zVmGeKqSZ3MAr
WS1LCp7GB/bfZ6wAE6n7V6y8Fz1Or/LZ2jgqmCLDNO1pPVMMKpx+yefpo93vGzGfB14NUdg2fmBM
Ltm0qMofC8879qY0IgOj2GrnFEZSL9gzdWt4i6Wlmf6xoh1ZnXgw9qH3YZI+aEUYzC9WLNqejuJe
SjFxJr061Sxad2lJGUQH7m+CaxtktU3V5x8F7W0JAgR8OxIKWWi56VMQXGzVfDTlnvgaP7OFilt6
96meUHhE/4vQqlfV7yKEAXUtLCJgNlMOQdvopT6KMz4sReD2y0diQMXF82KPD38535wou8bj5i6L
reibSY1PikJ4KKbSNoApccFzQjUangaVzbk07qjHLNTHvNXfBQYMrW2PgQG01xPJKoJMM2GbR5Ip
rn/M/Fk3r4CZad96S+OegGUPVNLNY9abTgxaqmDcNxQptmiIdgO+wcr2Hfh+vw7vKg0XtEWl/KSN
jzAWNwfJzr4ECGtfUCrY1muH8vOrdjuAE7UFI5wpQUO5BWGgs1MHgTVcRX6BB78tGcaC9zW4KZPB
sMUqIUaZbL+w2C1Zp0MW7tX523aG3V4YUm9VjPpfpxHd0akxpuC9tWX0OZRbFNRMHZbUbT1qFMWS
5qqNH8LALpCIkwL+cYHI8e8/h1QBXkgxBdiPFrWiM7PA8mE2GG48TZjG8OtM5TthbUeJhlITzkK2
R4pce3MIoylrDQh1Wv7lmxQJcfuzNvfoP5xwqT4VSEND/luesqJwkNLSD/PU+SVJzilhUlC5zhxI
LSVtIO6R9188zK9smA+MlQby8lhklm4s2aRzji9faU91qz5u1ijjkWiw4TrjgL4JR4duhbD6tQEM
ZP8ZBE+eAQc5o8AGI3wpDbD1cE8WHCImN21jDNco+xa4COOmSUwBST02qlSK/XyCZ1blBI6qadVk
KbTiFBNtEQwn8G8DXOzbVN2o+AKUCV2rzRS8g7HNymWHY/rfFlR464WBG7hs43xaLAdSj/ZUDhTs
Kx6it8FLz3zn2CcU/7s8hBlUsY5kyE2s1LqKZQy8/cbxrqE9pfjFPn1/4HQudSvmLJnCzixkAH/E
TRCxWAAIJKWx79BkxjoydEjiMmpaHsieYo1d47XkzaK3HZ1Lr9JNEre48zUKSEi8pZYAQ7ymxnnv
yqGNHtPZtO9YmOW/75rnqA9JW0SYaBnibuTphInsReUCD4ElNzsyLlIiyPErJArPMJpB+799fFZ3
yfU+l0a5FAGnZVVEKSmKNqmVAp1CVPCEnqBtIocfIEKB6MKSZK295TU7KrOGUyWIrxP/5qDnx3Ot
uU639TwnI2iKef+dxPliKhPS8so9zrZL9z+6hp+vkXE+O0pmlF8Xt2gGaA+1IKBxWRkz4oOGP1J5
tnHHj06FIdwiW0S9nscHSoeNbxswXadVCJiQ5hbRmV2hAKeR1ygMzUZuvxe3nCkVySBlLEBjuVbX
fBJvyfpJhLl/cSxM1n1D1i1HDKh1HMIPE4k5NkxxGo6IS6xRcNIGGkPnpZc0q2Z2BTiNWI8UhLdv
vxVpsznLscNE5E/Lo7zs2y+4LlsECp/awAAdiidVS/jpJL7SwADYs1YCeonso9OpC4NZP/L12U/v
90h0J+fBByFQwFT6BG8eDJHVvLwoYBH6lvck/CZ1Q8qM6esa1UOStRMdPB0iwYvngNpwnvkkUL0q
h6TdpFscb4G86y+7U9hYryTI+c/Jwb/gL65ScNNn9ju+TVsaT7ufdAszTgg5nrRof4iCpIdA+mI2
qNWj+tm/sJpzx4/cEMMw86sd+CTqcUEDKK4N4zsg329N4DLnzuftubNE+6hGSqzcJmyY0214+QQ4
jnRZjUi96tr8jb9iradYt8Zvl3LnASVFFuFe5fgLL12EeD5vCrdHGzIcL861j+InO1SZ0G4m+x/8
kDeDIJblvtpA2x6N/v71Xq84M3NwWNMpyA8VfJB1cLTI67I1JfmOmtSC6Gbpim+XlIF7eeyV1TyN
DXSil42opmv7Kj3DGUTw9TZTN73a3mDWo0M8Fck+IsrZh9p0FtAzJlPFzLRq2bCRpnHcBlQldhAV
tD5hcXyUrdEUAFokaIEbSyJvAnOiGa2a0tzEFAF5LrOhqWIz62CgrMVS348FGeK885xsWzxNSCco
79EDIJKiAbbaYLA5lAM4QzZdhwgahzhacrYUgeOehs769XLco255Jphq+0HRwmpSdF9eWAH3xkmI
lkxoYVacLOK9+Q7x9fKHzftCbL1tfNo70yeoxEY4O369P/BRA2HPSM2XRm1ImrohPlBwsVCiTTgi
KfVOwlfxPn5vAAvQ32W0gaFh3gst4Tr1geCCGUantwK/DNbc61dRHThe
`protect end_protected
