-- (C) 2001-2016 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
qfta9Sqyadhusqpa70HkJx+nxIOgGd2rJdslfZw12f3Jt85KBU345yxDB0HSiYmaqMZ6MO9pxynJ
qAOZ02JpwerzGDekjK/hs/5JJ+y5rVdQH+ifroTjxadJGoy145FD6A+RBSiBwmDRFZFml+ns2QIX
huWyOKrbeBx03d5X6phKcSBiBSx7f16x2Z/zgY4FFIInAWJikOxX/1ybhAZg1VTaz7fIVrmAtmFZ
7WjwdzMW4jaubtSQfVU5Kgel3QeNeXBwrhYiABb5VMvx6nQN+u79khZHycxTyJeo5gaHL0aQkxjS
gTiObLecMvJauDCgWCQdbnGHjRv6yLrPljkwtA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 2544)
`protect data_block
AbJ1v7W1SOJjVR3rYCUQ+Ukg5dDnnsLqYG0W5Szud80WKB+V4ZfQAfAu4ZcGLrDgLd8t3zvYbxwz
5S/9I/AwQYkxVF5rkoBPrMOCiy2zgS4otr3SP8pMpb+/pdnC4ssje2Ak0Algltbav+IgzQKZaSe8
QXvr2Jol3uLbHDkVC2FJA9j6SQlqk1S2bWyLcf8kEP1VozRO4WYUpfzcd2GbeWqalSY7hoPudjpO
9Ny0RQkaNsE/I9I6bg0y01XKObN4G1qs8Ri9Z9Iwh8JCoJ5A/11bRonxkJ2yJJTUxUZfEAjj4LcJ
W0+GUM44iLPy/Z6BZ8ijXNb+XfLrFcyxjFZUdq0CmQ8hBzHlSiI4k065clLnw5b+37tnPH2FX49C
Gi+gfZsjTwwaWjj3HKQKPInCdZOdoAof7BKd/D71b5DVaKy9wcuCN0yR8rF/rcN/1wuyaNzYlAfM
2gDeAiJeBRw5CcruhY3vuPn0wNIMJhVzqi5PecQJf1foP9HxxdbzigNV3GFvbXIp+71xKCmZzVUx
EWonVHLcTexfda9V2T6iMCx4P3Ye8WfrZy+9uF2R1NLk+FH0N1cHupAmxAUtKKaAkYb4PUsWS7nG
wYY4Bqs0YHqVwf9N60jfW/HPDUJRWFisIT7LeLOCiBrSph5faCoatn54u/D04pLwpMazV5STynvR
bcHQdEtvyTMVgYX/dBy8QE4bJ8SH4xWBRhQlAajzPwYqqBQzzgCMtqG53ID4nVfrCVcWkwbGBccE
Zkz+P0XYjD52t7SZf3KQpG+tsBJWS23uZv1MvBozI6pJFT7HgdbR0H7kFtsQoBlD5dFsCKpW2Rmf
JLZ01+w2My6cpkUiT7b8NL4ayNcJnM2VzwoLy8Cf+SonABihrtG3xrXzfN9wrdinLjRDoB7LfZOO
A0MSOwbKHFDBynf2+fFsMbwPzn16ua35fazMJJtEJYUdW0LPw0Dpu0t+/ObeWbMT5vk+CtP840b7
NXj3Jbwunm6oz6sZP5rSLmcvCSJqC2v1vj3rDsezPwTKavodRF+3w6mbsgoaYfC1Sje/1SGTSCON
tebV3hoD+kB9DWbWpAdt5PXLnOqBmsjLPEkhO2AvmZDi64tLsyNWFatDL0jpkP4F+AkkXoPOLFXK
3IJnanv6bmSMT2SAmLHlfFFuVfqVprQgKxlgwZjgmvvDNmfLlAQpD4q5tO6Zfv8qHmic4r9wsbUl
65bu5S9XfW5S9waMnzunKfcd51pxYORIzr+M3atx/B6CwOhS+MxkoukKAntfKhrCgSdQ4GaMTJHY
oqk/bzeBhGpKzeGiqNZThCvACDw9Savj8OzaAeRRoWnEAi2HybvBV/0pZQLvgkUbwX1SBuzj+zWB
Fg+52x074E7/x7qKqOmNKs5q4bZYWmgExtoB0QSgUu8Vwbqdwi/0G+hTfNfdYg18wufSf5gPzMbp
8s9VuJCbBTZ1V/v4Hkb4XoKmcZ5M/PLkBZ9jrCsfG4jNtAXz8bmWGIDZuWrEcHvIpyxwnENmzwLu
0bj+r/MIb8kWbnRhmjUHmDNnXart1sn0riSCGCqHO3mq8A80y3TRzKS/AoqwsWsKLKImdFsLZjF+
vZ1qCBFQ6cP0rkbRYPLYEsIuoSmX/MrhMukYF8+NPUWqDbYdkFqmJUIMi+IWQ4wNGB/08kWrztMf
+ixOv52HHd3vseXUrcVsURe+ak3uCyLIsOfeHNVIIgs47f1fRfT83alLIG5Osx93gKA03He7dh2o
ShfU4ZVZVhsmH8abCaakbqMpxag7dIm61O5G0mLPoZkcEdbBTpqtFzXqnu97DljDApukXISreERl
kfu1aOfDaC22OTVRL3Hf7PhXfbb4KMq/8I8mBjgty7Uk3zTgfBUXaxwN5kWCsg7nh68CfKKDjY/+
eR6U4ruvxv88eOWPwldqL9Fex/QWbqzKZWigKg9tAbRpNKkwgFZZFYAMZTGbkEa9GUdmya2KxSz7
qqPA3/nMl0AHK4+zv/cGWefdBtnDPIlI0xaJRlocOEP87l7y3rojXoSaYZoEQVgRXX8T8dFT96Ue
s65uAchpVjjE8ybXHulXLDJ6LZQJ48sCLttAve1V2FjKBgap4au7hDM5g5ImTYF3naOqpRdyR1Ib
JWb1eUmh9GSbrsWULKq0Kc0HgxRLAW/xIUSHXGTlO1diWhunX1K/lDF7PvhrXR6OUK+euy9+sFWA
J44C+2r+RRiiF6H/x0wRey/cNcgGizLq4hyNjckl8Yp7iwyo9IQbKYeo70wXInAoZHfyMl99IKdo
vxehXPtCl0mbjRIIftsHhchjysaH6ULJcz5c17JRv9ZbcDZF6k0xnNcCWHGp7SrJNBd4NbMuiSEd
s/ISdnqg0HlC2XQk881rR6a4D4XkjwwMzDUh5siLk9caqhIWNTO4KcTlGbSc7rVke21jyOwaoC/n
OwhESiQdYtwx0+/KGhy41uX7HfYfigdvYQ5UgGrht5xiknXogFq1nk2hGQrB6Hudoa8qIEniGwd+
G4GzUwRzi0GuStWljQPmWyioih2quvKD+IW1YQjL8tOkygPufK3PgDapwPPQjIVvQRuv4w25A0KW
DcJc42bPqoJVcucN83yh3VtOtkPq6Bl6hqWKni5zn+Oe+Tz5e9L2CU6FexdOl42kOEMrwwYJJocR
Kz5/kMseknWoBKkQvbC90mjys8enxFPNr4PB2ezS3kGP0lDE9N1bKIDgYYbWFXJLTnnJMfsm20Kl
hkvMw5g1QcP6k+jrhFo3mGL8k2AsN+2zIJtQ6luw6Zj8gwskFZVkphtwwK31pWfL/nDJjaQPOJyd
zgIRCwWvsWzfP7DCLcRIAKYxwpryUEGGbtgb5HRN6kpU3kSvsyxCyHLRjS8CZJeS4Ki6bZMi2tr3
DXATz8OJAWM1aJV2bqDi2golXbDN3KeJ9YZRilLzxyt5nTkLV64DhxhU9dRXqHur/LV/DV85ncYN
fbEeyhtkr9HXtJP/NYAmMgW28H9uWftXp3LdEXaAvxDt0+660Jx7Tedib7JQeUeZxKYb769bHsIP
faotDNsuALAOVTI3lQwZik8lueN7YsQgJwk3NmRK0zZqiu828LYjrU7lSt6MWkqMA5LvWmukaGPB
LearlC8LxcfK+SFIfjxfdh+vy+LgNaQva4+beRbOwoZcMa6udJenzQfLRUNdGnR6W1d7NuvLfK3V
NNmca5tLlJF19bS0IJVX6WvOPEyGIWgFvMKaGQZSzrw2VgeW2Z6cpxjmscZg5jWqwu1JIgVvCs8D
VM5Pth8fG7C84aEMQPnNgC55G3xlMEMFFOGDRR9P56tzLUfB9Pb7xLZQ5Ps9xwOBU772Ofw9rgfS
wV0K97N/a8ZZE14sIcrjiU+r+byR0Sv7Jtrc21vazGmk6Thd
`protect end_protected
