// (C) 2001-2016 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
J0hOFxRc9DPwgx4NXb4fpNmf5X9Iyuyse/ofUPLruGXsL6Q3kllNvtcUHIJVwlo269UV2RqUAOth
bacs1aOWe3f0JeLck/N91GfHIvF9iL8/wbTmWN4zhEJzqiv672MQUEecsQGrUCiAh9ygGmlT870v
xa98JUKF1xMJtPu5an0qUbX83z2J943tJ0fL/KOQAwNjhEbDf28faEcTttjdwivS88BXE8rSje6n
gPGy0wx/Kj/8ASPeiTDeGGtHmAh2xzOniQpyMItu2393VgnAT7FDNXWwqIMUs9uH21HLlLTZMM+r
9ZtIz1dPMd+wDEDnuhw4/hbOdP8uOh3JlIpV3Q==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 3936)
RMXlE935MZfq+97Ssj3ePGO5q3ifErIV2ELiczCLEePWNKUFbeLe0mmGHhqhobWHDhhGriT7OKEZ
+Lr3MmjCHUyE+QKlNLLyW8B0BrveA8Uf6v+NpE87F+Kzs+frCoStMOrKjIptpkn/cKcPmM6Qk9c7
EHXUfOBPABJdSChXwAuVZFS1vBwoIsns667PuNoQWEezK8RuTHbqCd5VVHDbq32Jzhz3YQgEuKcH
190LnXoXLYbxM6zPPCbCrr6GzxiZ1WCX8i0Vy8XSmoP3V027Oe+n0x+4uEwFVMLCIRZp+lUhqD5E
VuMbzMaehcM8WFTCUoqUpGhOSh63YyN1ar32hzOThgKC0knclJUUjMWCvocY9XaLgNH96RAlaPlB
TSvDAsdubhCEwR1KhXNRdcSWb1m5/FRI+MQqVNoklTMZQ5QdJlT5d+MRjWU0s29dvUuPMBwecuMz
NF96E+KNa/AhVwhXpzWLXSIFA/rHXC60fvvAyMF+M51cNJjxMDXJl7MZRNkCpIW8qAl7ydsvvaKi
uJFMM6t7+0V9VsUcsyIFl7jvbgzDrcGjjOVZE4IL1jYwQtYgKLrv2hU+YH7FQvHi+6FD++IEpDQo
2rvmfGPVIPd9uJ9p/WhgGalm9fL5U4kFHfhqiXy0ZY03QLF7QcpPlRSX0TBtfTpu0l1Vm4r38FhN
8Y6wORmsPkcyvVGc0djoJCbXBtIX+UkJzUntGoOqwc9coUH0IRUOIFWSrqqX04YWsbQyzaUkpEcW
E1/+pj3Orggyc8Ou+raPVy5srEsknT1o8pHTq3v5fBF5cXoWOdEd4fBFknqi4keBn4AzZ/KMH9jY
dm1sPPuxNp9k22snTBBcsz3Airo+pfUlHSxVgnsrXRNt2dk+9MLaRhyASw9iRt2wGXFXbwOgr4ww
OnB49mqLRBb4oKp77IOl8w9KNiDDX33+8ttoZk5XlYI5A1LETbvHn4+3NCLuclBe1HTg0USgqtFQ
nm6s9q2R5QQHQNrZ5pvdJP/hwxeS+I1f/sqgmq+x88ZTU12qa8GKZeQkjtg5WBoTnw/mvGpuu8P8
dfO4j9Bx6/FXcPwKcuznLWwdpR3fjJvvLmVFvFyxNZi9SMnQY7Bi+98dJaRvO/Dx5pd+FaddvUf3
yjGi4KyKTyQ9BkWhqXkpHs3R0T4yqRgm2lYp9kqXEeQRVyqCnVyW0oYRq0HWwrBY1a7t8eSPlnGD
SfctzOCmFeU+x9hEm+3pYAUpuWt8/AZgqUd6AHlMO2Ya6eFzGATpyfjO5hGAYawz7KIfJyuW2TT3
IG++9VjIP4w1DEJ6Xj9fti0TnAbI/rFkmvUOS+Ws8n7nYlLKyKQPZxFYyHwFuMRpGqYfYgguPJDf
ye09009mZ5DJkZZBOO6TkNx9LuGNInggmUgKJZzoTiFnOOYgX1uKqxnTgxpXjB1Y6nnUth8AChsa
YDZWQWbX5Lztd+65FDV6xgq2oaFqCx79lgIsN1NL5/RbPmYhsu6uNmmZbZKuuyfUzzlrCvd5jodG
fMqqvmkXQFGnuiwcOMOJ3dxG0+c9aaAUkEaZeFPU3x9iL1tpsWSzLXG5eQF8BKiDW4EmZ/2iIN/D
8BynWkxZkgVkwDVfysstfMDO786kffYMimlOX1thtXkNqev+Qg1hEke+NZ64nwMbbc5gbGjbBfwt
2iyAbolChA1UR6CoamPKwv2C2DUvkOIcgqPCwHG3Oz8TdFCC8i2MrV+RePGnR/akUMrN3AYz82Ac
JafS8jLf95uaIWm3L0JJnrYwajJgwcvK5lArRYzoK6ZXlm+k1JLapEHn/SbU4qk+nRbR69oMmag8
f6A+a4a2h73Wnbs23WZbCzG0v0sPGN01Qc7vMk1W7ysn3EDgKLo/o92Yx3gohVvuDBnQ2cRMk89W
SBUXSjSxCmc0h6JFmqOUo4GI83HXJHNwbpWX3HBa62MjtHa17BbQH0GgpENSYploWoAomlGj7Lr+
ay72a/rlADoGTJzogVhNbL61j5WyOLxv4hdgMNVZue3xbOfXmTP66sTlBHiDn2WUMT2R6kL1cx5D
PyRZIL0Jm3MERF/w8JqMdEj1OrOvFKRlITk8WfCUnWW5Yin6MkpKOy0bSw/Hke1E17jlijSTJlB+
rSRly+/7cxGRu8DzTM0QHlAPnTehlDuxRys5IYx7rj6NcXjy2HMzEIQRPVXyNP+/obghokKqhhy8
p8nXF92M5Xkj9CmbpKUuVDTQnGCJBwHOz3qERheemGs1irRX370jijcF6wO46JQAQCsCNzTf3Lm1
KD2G1oFKCsXGWS/qk05qSdM6NGzVXaKkra2xNpCqTTG8WndLb+2HfWH7sGQ2u3rihjW+SaiYNr3o
i2URaEIH+hyP9mRP/aprqukxlXrFk+nRj7PAMRVnN7pDO8pn/hv+d38ry891xI7+qESNfDKDoaL7
Ge+9BHQPEwpf3uFzyQ2YwhN2Y/e31SalZ0+gvqvNjTb3TDYeh/Po63zZewpxcjPlljjn7QBf2jdp
PpQqrwXX11RIja03GcM4U5mVm8af9+6w+ZbOqyvlDzB1sIug4Zz1eDgOU/JEPHnzqRBOk6L5cNLh
jVDGsnYfBrlCLF7lXRN0hYbYTYgaBgKNgHOrMWDKLUXwhOpURZjRZxv2nSIc/IpyRAXhk6Aen0MU
hSCnbovNy5Wy4HNzE4fbzGQbDLI6MCQRnTvuSUEhEdmIGKs+i0ueluouxbc7tA3WYbc24WEIQzLa
KFNGDPifwjiVsaschiXrzKA7fRcQVihaKrv3Jez0vRlJRITJOYH8K+clXoEoUqwRXh5U2Xt7gLhR
PhvQpOtKkMFWd2Kzm5sY20L1avRSIK5fEfa91IUNzS2fZ6mArvjucXo0MSg6WscrNOeOT3yIfzgu
45hmKpZM0jdVXMWuV0ev63JwWEwTyAnlQ5yWJzmMoYtxvpGQMgOvBrQi5dnEDvgHlKJA+4pRIMqX
AM45GVcElkHGPtw7lpHL1DJqn+9hfrXWcmNUpEmck6xjcwOOzKDiPhqu8ZhXG2TFeCY2YNSEyAcE
lqDytosfCB3/yMUkMq1WrZxBLTcFzGIXvQGXn/O0tLwm+jDuKGSht/fbsd2x738GKXyX7I9htRYp
jhh4SC1H/v5JqPMt/PQXykyf4d2n83fwWA9XGxo7EKQpGZL+PH0dJRU92ysEuKedehOfCbJIObA0
VkMdvGa7yk/KuFE1NWZZO5XzhAdkzm13jHYBf47yybn2e5vzw3Uf18BqUhTvPSoZi9DQG5Rn2NRb
lp/bdt4gctuqR16SkeBaHJAH+wPzrq7CZ4Wnikn1/vcGho2gfiajNG9x0NSjn/V54Hri5NtshbXO
ueoravHEcmDODoEoflC46EyTbkdxZIiz+HfVNgREC55y2dvo1pFZlVnLCGjg4U9W8RFStwZHFfvY
JCckvBBCXJot193bodPn4APmWW/BOPgPZMuA8utfm24rKjSkKau7Wug+QZmROqR4g54Ay7tNMPLs
phI3my3wDQB/Pf2CccDf9QhOtOVsVWITsU+TR0R1n1e9N1mnSn5rAWZjkhcQA//LL7P/XqETbDfc
IXnRN+hVknxBN6CFvNdrIcNb3SQuRPzhRq8LmTajmtu+mBkOs064XI9xIpImh8SjeYo77C5uVmJ4
oy3iG9MKlJiw2+R/MnKUjv/ZUxzaDYzYEK2V+5nHo+shT3qHx+mpgVFERv4e3ILr3BaVN/827da5
VP6b/Ky7XSimAX8T6T4EJGFA6WJTPpXPC4m0TjumoPuRI5z2hcL6T/YOaUzAlEYjwhnH1DpUnMKn
UmXHilLZNGesbLwLgm9uTNgdjCoIc6Gvi2xjSAPQ19XdkdGNmMfW21lyM+AgqMFm3NU8zVB/+EbO
wXxkovvcwHq9ld8oAl2ychlhVub6tqW66Gp4VlIokLRoDILyN+v6um6qSXzv1RCMtfqVXHafuU9j
7BWA374/WCncQ4C4i76pVHiI5/0heRQEeQEiUh87wg45nWTDCmV0LmyVhmI/MPIfGEfxDP6qpz7c
QSmQwkNs5u8zWhnTEKLq7htvXGkMZY3LRa9dddrakHFTiNJj7yKCz8GPUGlJi7R+xShrxFYhAFGX
JJdVVSJrQbREC+4d7pyFXK7YX4FSuFD+eUPxfeHz2BWu5YcJOFdEU7Aa0+wdeUjwk765eI54fm4E
QbLJTOjH911hJ86Rd9sDsSZOfa3OUyWRTX/Cjh9alfpeXWXDrQjD8I1EbHNFqKW9aCIwLodCPgc4
w0lsSCDVjQuSlRhqhg+Gm4f6eX/p7CCHYVaZ/J2CqtdKPsvx4Aoj8z5mIDmfl71SQS/737sq4TIM
Z6E57MbDuN0++QkMa+qs3ARQPtRf2mH4iE1+I1U5EwgqKhUM2+32BW5PsgERUrTTFQexsjqRyxgu
PEHP0IPt6od75UHVSSk1U8EXJe/D4ZrlbCR8UZDCQk/LELmV8dvo2kHC8lRmCxPGCTFGXrkRHh71
BNZ/LKlONVCStKx8mZYFVibzI0QN/kf+DqoZk/yRXmlx5ST2XSUzPXqhKvaNjFcBKjgZl+5jdvMK
dVi29N+Y2j8Q4vLXJXXRkjwN+O7e2VhihCKUJNg9q24Mx96YaZgesr89aDmndKfm7Lf0gEuSNOFL
WeMJi7dO10QUzJ/569kys9gAccdZdSpWwDXj9jfh6jn5NEohP/2UQees2TMlx4ijTdQzNd+SAT13
vAQikc2TYQmzZzoMjQlvqSkq3mkgBzHlVr40MxCM8mrFU1h2beymLNhYm3V2n5uiEnNjfSVt/qIY
D+GBKs4gi5Ix24XoXsmmi6MYOOUtho8oD1oOnFmgUxUX4+6TE8KP0WPiZwQL/bmrvDUMhhvMvzRR
1dVI1/ZvoIQZRgmQBelg/8hzNJCl/+WfE+w7Lqzp11ZoXK9KMiKwDUTqyyj3ASSwFqEireP9ihJb
HPI9sppQcFu7rfjB/k+1vwfQy0s4wABX5J1EEMZh7nvbAoS14lA6I8ufkeXspLEjz51G318v1bzO
CX2uuRsiUUJRNjlinoDmeu614KuUlxiPnYSlaGLbU53MqMALnLzvA8FMG9rdQHTD3kpiZumHcCeN
oIfdCv38iZfIn9sHGlRbDjyIn8ZJWuvXu2hjrzHIfdeewLCXFLzXRCM5hl873MZ+cTNS6Dz3FomM
UZ48enDeDB34jYzl4Cck5xhRYKDpg3LoLp6PSYlvr/+VWDIEhFNG/8ebWWKHr1s3nndJFfOMMTP0
GZwD
`pragma protect end_protected
