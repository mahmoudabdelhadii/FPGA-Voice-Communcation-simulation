-- (C) 2001-2016 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
nuVPmKipJghuau9iqjIzj4z2TkpW0KYxqVTX7BxAFJl33S4v3vLB6O83bF9K/FO0h8bp/CAvJWpN
usAfjoLMiRy4ZQ1vRtWqep28MxDx0Yz5shVdEZDOvJs+zjcG+z2oBmQ3yPxDAqU77+izIdDDCNrD
4ikT6hUT1i5h99NJZ4R3peqOj42RV1Gl8skKWQKWCUr918CnlQK+D3RTT8fva+pbBfFERbSHm9B6
gsN3Gdjtdbl409Q8Gz/MgDLTKmgCF4i470nxYozUPYdfFB4pK3ll0tdhjcLcu9uwIc90Hu2oaDoj
m2KkUh0a5YpKoTjtm6OP+75QGP045vgGQG8b/g==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 12464)
`protect data_block
xzcucV8Tda2dDKl2WY2Pbm6qyfF+nmwPsChIX5GsrQYu0sB8wSLwLzLIi7iyWRtzdVMTunai1JkV
5ZrJG6IwdsdtGwfOXNvQq1A8TZpCo3d0MlzuppwC6FCMbg8xatXUTJacHqwFfGfv76IHs2vkUnsA
xBI5ud1jHeK+Imb45W/0QfXF2rNVuWk1f4/p8qWTIlh5e1BgBpzRATYbTI0gQ65WLvAGhqLFr6mT
ib7QygFI8ED3HzSmKcl+ZfK31r8xvavqui5Y6w0CElU7J2iQTSdTkISY+srbKcgJT2UwEf0uvdMZ
S1H0Ssg6DHBDFfBSieWXDelCuMetmgNX+XSlq/z9VfIsF9yfj0qwqYRgeoW3Ygh1JZD7/upjz6XU
Agh1txrts9H4+Eszzus+OCDeOx9e5QugKJ9uXTq/ErJaC68+Lg4utqPQCAKVKkhASdap7PCPEwy6
yHzFgJ+NMPaNBg3PP4nTM0IL3MPpWriAyurAjqKMrncqlAZ+dUpM0EiBRfWPRPEEo8djDf8vQ/X2
Lrute1SqHObdx6rcS0dh7+gnFR5wOGD1HAWCySYvLwsHx0urzthS8vp2WhdBUojunzD3QC0K/gFm
Ops14Y4Q2WbrD5iuud4bTJpo6VW3ZdNO0cEaxj/JfbXUjWPgL7ofSfdgIZj7IavAr5b98dGec/GZ
BYQFNlDDm1iFrWsbG5dHoLHO362ZESVCfRyy9EHMLVFP3wM5pcVE/Ihd4QkbcmDN+w65UGwDPp3G
fkd/SKaYl9Z65ft/QJx/y920Bryd8IfajVPJmOclLwyvEQRTFFRFUD6EE5W/+1Z5MjlRkQ/G/0V1
zaSwxkHJsJRE7eSph9b/tS2DjOhJXZCicp2v5x9PhbUjkbQZeJd2++5I1TgdNjLlgp9h2Vf7hwzZ
PEuY+lDNSbE/fOhhRF/nN6g+VR49fr29J7c/F75+Fjs/JaHdDe1n6O/C0B1MoqEE8ALxnhhKRimt
6kTVGNSKCtgpkZpdYuZZNedrvtDWxyMD2eHSTqDkl3DLEmcCFJF/DdT+2DDCfJ3cP7OCFJqq2uRy
arjN/OVFnFO6K4cEHCS7tGYBnfDtn4usWTOAqiJaBZLXlYVrZ+Aze+7ACKS6J1xVP6yEM6VQbyVu
z+eDXCTHRk0zJobNEmadWh4bSmBVLiDXHG03pV/K4ihG9bvopiKX6DyQh4FB8ryVVd0bj+UiMCkU
iTSMwaXgWGxhv2HPZXKoBq0Ds8mlmBZVbsLKwBVrrDbCw/8hE8msG4ibjwptlFJ1XfewYb8vlpTd
j1O3E2FZxaUejxVmJakbiC+jO8WlaC3/OCFxz+t3kyKbVYimdNQ0KwN8FknK1GNxORXZd4Pxrr5b
D13nhXBP1pf8wu1H6+NlL7CFx9b6n0sGKfrwRPSDrN2BdovqtIirg0Cx9hwf4hxBnASgJcEbmnKl
TWS1I3DjSH2aA/c575DiMUizYC0FfkW94rtTjmgxp5cKRhAYJ8CS/2vF3v9z/bczsuAXwWT55fY/
n8Gb8matqK8I3mMrZ13pX83NQPr8k1ruB6bVOvvw+gClun+OCb1n8Eaw1UNG7LfQUUkzU/rML8IM
PCcPWKTmBo/459hFmE13zdXpmloNRTQP/wWCH8ZikQdXU7W00JXDPtjhadiBp23VXWABjeg0mPck
mft8I6zQum+9djMRns5tbTjlritG67Ykfe5cktCnNIXUoaZ/fs/IPQ/d65G7NGPHmBcMp+qwixnC
V3IvEZLwtEq8q73G/HVUTNbfq7HMCD3G9ZY+CS5Fy4+MJnnI8LjxJpjtHFQmZvKKR4RQqwVyWudz
W9uphoQRWXfh+mk0I4m6sIK6yVnqmlKmskfz0UEaJNxe7FYiYXY9iiKEqX1T2EgKilegMf37VVvN
jC/N3w7PeK0dZwT9wZOiDGFG1TMLVVy+ndQxWF8tyqDmbQbzE3eQ9IHxtF5zUknvahkaYG5K0SLE
7Vfe2jd6V+z+V+9D8+LZzCBoR29WGrwI0y5ijndOGlUd5ky2ieukBOF7/9qMFK9PM4fgpMEWQf4p
T2I3V2mxX7vPLiZi31jxWuqCmWXFoUjt7FEKEq82wj7nnZcT6cz4R2D2AcOEB3l5YCGhH8z07VJN
WFWBx+HjA7NkZMgtyt4pK45ztAEGQUFkbpSir0HF2zEk6AnkNnBULD95DgoHq8llo0ZXQcO+jYp2
IvyWiSloa2FDLXXu1xkixm8BWOCr4QX80ZyQaF30iQ5SaWmQsRHJ2cWaI64XbCa8CdyjQuyPmNWy
yZkmwZiwU4A6a6M64XN77T+yP51hLkZNYDqZFQmHf+SfqVzWVE8CzLTNZspYkL4ppfQfYvIDZut3
L1pk7owteiEyAyp8N2Ge5WzWD7uLgf058Gt0xTkmGWaCceibMo29HH8kSaelM3o805oD8r/hGtMz
O2plAPcMfFGKTialzTG61b9nQ8du+toKojFwLAfJQLYPYOry2mr4i5GT4Dd+zqwUjjOcp986tGKT
zRZvefskZPdujzgBfOIKl9TFzXNBuaMH38zB9/kTULNcwcytQkTjON67oszxp+9sE+QqCLhuzhaN
ywrxqBEpkIafcinbXdg7pE5GVUVhxdSOuKvcYLoEBKuW4LkBgMhkEKkbo8Eh6+S2dkIKagrfEkeI
IUy9UnOzt6WCi2JLBKdft0x1eIVAZsFsI+6GvsVS/8846XbzM7fNDEYRyaFlatdfBuraZO4LW6kg
4t5egthMIoJGnHygKsnBZdHhFVMMGxnq3Q5Rqh9OpiBZiF+XSadpoq4eJc9q/8RrrHn16gCQePKr
2V49xRlc7HS3b22Qaojm5TaeM/GM8LxR591DdktVovcUrET8TQ3ENqB8tX1K87Ug32DK8Qs44WrI
mYCoXI0LEXawELZklxBduJJa+0Y2iRweS+XgClEguxOcYUky3gcbkmn9nrA7GHGaEyzxdfBDLQhv
fN0ldxMDlPMuNblu/WcYzi4ispaTyOgn2zIIQpHXHIrKQbo9mT1QthHFFlXv83TgtF3ZbUReiM7S
cBZ7FEty6vVmfAGWJDA7KjMPBOj4PzTfBDARJNYtPoy7GqartgMJ/xDQOFe1SV3cYha0LgwJiTZw
8QNLv4Swelzbz6knVDVN4465f0rqiM4P8h5uDc6jyRtcS+fODMER4oB8XjJTHZGKuURjj4pBul+5
lg2PQSDs90tmx6+B/ImxjE3bCIznRNZUlBl4wtio6Xx8+45ESp2ylZQEShkI36/4EDk6qJ6rAtNo
x0qKRlFXECvw/IP0iiyTtjCBftu5ohGICcDC9ypyxPYuDKykys8HCkmLlZnyTb2R09RIjoNry3He
LZA07Joru8T51UgY0VHGS7BPOECThT0AjjCTXZPDJ4ek5NVXk5aLw7LM5OjaKY30dcSZ//9iDdQf
XRSiJz14N0TttZV3M7jma4k9NWYe2mA9NvxTXGyxOddjTDUW+1obM9Dn4aOto/cAalF36/7Li5fo
EEq8p8CzUBU4ARLf7dGEFGusmTcmkeGBY/bSwOKeA/sYfWIxywTbrZFGvw4xS+Eo9Hed4cftAtV+
6amAQ/g/B6FrrB9NBnOFgYxifUxR3czuCd4yu21UtlvkGaB0wGduqDSzJWQmLzO8DmhKeNSxSa/m
6CPg/g6IYiosfDKX1enVlQYjX2PBK7oB12GTk97QNp1TqJRAVy5XKFO6Gex28xEbrNWRUGnfwtOJ
LbPbeWYa2McmD8O885Nnn1pzDm5fHxcJW9V+8K5cikuZumUEHcRxI81oESJ6hROmHjhoZMY6y/Bk
4DdG96t8D0BZxExJy+Y+aIjZE/xAwacBtg+N3yzlZSlxjokphywlaXSGFoRDCHweql9wH//N3X91
jAUo1h8xe+gHAowxL9JKnKwbgeET//nhbtmWn/r7GCI7HjB0irlAESn31rbomB/yhmk++D5bThmh
mnLu7nifqIgH6TvDxTPELeQzAR8sp8Xy9K01jfb9WI4b9Yh7pnzIaBg/hwY7jqYEIZRM8tiKNGHj
8TRIeIQqJoCUW4t3d2QfeJOJisGNwRV6+aBxeTgaidJl/+aFJCrHloRAlRs1DOkX4F9dG2F2GS+b
3Lt+Nd53cVEnqkY82Nk0fInkRIkXbh//znNPPjeOaOISEAHSXYhbOr50smeCCL0T/BkYe4g8PsOl
lLs81ZYlMDyOO4uxd6m4tOd0+sNBg9g4H84+j+BZUy/SPhG2unZ8R8xTLFyl9aTzGZlJsvL3EFYO
x07wV53GVPcSJIhFrr8yrnIIsCWgeNt1QHHJT0//P62t3Hf8aMpSI2B1x8vxfHS+PWVGmHXLmyvN
m/iD9NzF5I0ZYbWV02OCc8rc3g0rhzcH+3oGheQS6wGwRXymPteq7thnLbhvJomHDB7AJtggHzM1
Sp9k9Wqb10WkQXFN3gNLbUz6UwUyy53/TEGHKig9MrnvyV4BFsU+W9BVisdh8KojhXLwD11G8I3H
glxscRMlJIlkXWpiDjrWIwrcsI+Wag4+8xl86LEaFRJGvT+IowJTfmFkeUnaWgFiI9HX+kol6P5O
4ygQMRUcEmBWg9YuLio+SPUH18I9zCwNq4GmCeF2g0myVFhLSUbv7dF8skPCjfhSQ0+gKNy8MZ6+
w2Ei7ghtEU8wqDoK3wFqw8atUfspMJSi2CM704rZrDY7fCxvVe6If2NYAz16QUJ1CS+qwWzdbEm1
nd6krPWUfZSWVbhONyJ+w+USqeit2st1NgXtAkMqX3XUzjymN7Cn4hTg5JTzlvGuel8ppmQJhYyS
Y2qIL7W2nJVcfDk8fbhNZeNYyb9fMis3NT2TrsQ3bsMuYaVc0rchjbzsoMIaOggLTjq/LSB/6hXX
w135D8lJxpwdBgs0ho+hsbVKQPfe4Kf4GaV7r6t9z3AVYmQbStX36326qC669fDQajYRe7IyyBPJ
FTIJhuKmGqK+VXx3m75yg9Ho171Ofq0maKAdfGcbI3oT9KSoGu1xIveX1gGrJKSIRolDNcIO29KY
wuB7DrMNPDsE5m854kGf3UNhY0NgYpeg4lYnL35fDtPr0bpEfdHY3XHKT8bd62NITLm1vxipqpFm
KD4ASMbaBUlBkjTL0f+pl4OhYDUwvXBmuZJYb2t7XFymlHwdMazRGa3Qokw/aSg4TEtbCxdxemBU
n5TpH/fn3OTgpeuXSxF2aUpTpV18WriNxGjmVJt5M4fRvM46SYBL/2ehffm8V+DNVCKxXFcJevMX
RBjQ/+zJBM4CXWRsCdvoaatJRZmMLX4un487hL4qp85QkH3NRPJnafWN71B8F3Lfi3ogIi7d/Ixz
fbdpC6KWfHUxg0H/LfGnPCkFV23/saMnqBI+TYNOG+w4kGtsLePVhWKgRGuD1KswBXeRogP8Oljr
WNsldGob4TZFy9hQZ+8cR5advT/b+KelDg5Wh9MQy2DEjztN0n0Qr+MTXS2/3IXr3pNlKjaG56YY
WpbgsoBncOeBQOmSvnI+GtNHhdCTH29xoggvIAS9/HL+tb/VblUYtaFzmo7MU9iInLsSTidx/cO3
8CnmLVAXHyc7hx7Xlct834peYMWUAKDwOhdCsqzm6bF845rKovTN8AliLRbS2A/HuETpSMJMjOqu
qMn8ZA2iwVdAI/IclU8nUN5i1wAjQglNj5vvJBiwke9gBjvvR866SKZ2Lcz/vkM8R6+7eqEDeTjM
h3qjqlul0ZrAUSJQVWXn1HY+leUJOBw9DSQ7aeiK7ursjzyfY7wEabYT0AA+eb/zj1YgAemy3E8v
OLqIivBkjXXGTuEniPOjABqmwRtUGpfejVwfj4C9AK+0oiRwIsfi5cw09RJyZkG11BkYmovD6Lwm
Zuc0Vy9tzMsntcp5zz+BfiAK4Wq4GEdzgCur4Kq78CmSv22y1Smdo0jaL8P3kbjUkFn/RKNFHVdc
h/Xa8qHvsNk+97k2xJMTybPLIodirHesYXn9b0YYKwmRZLVbxOtOcoTK9Cfo7w/b0RsH64XEQU92
YJhMNtqdfx3HwgfZy+D6+Dewj8V37apO9+72FTLmgEFYZVblXfFKoKzdkrU42tQE1aA5MRlZpa+U
2CFNCvmfLb9rwHSHc6LIL54MiGs/PmsIUtOX8c5KOYxKRvmODibEA526ekGlQmsAExVhKapUA86H
6M/kw4Hc8YBO3ERfDUkZokb9BwgxG6+kjqmH9TTdZSAZDEX4XEgnhW7cdMTvzosr9NhvbXNGQxFV
ERDF0wlt8dB00JkuadikzNtiqD7ocwmfoHFoRgwpmSP9tm2H0KI2/0yfPqE3j8K0J7xEdJauIYAA
n4KYjaHid5/Q5CQ/Pv8XVKrnnE82/uybGS3QxPyvuVcrDI6LDrbdgeyKTdMuGMPB2kuFebs5ctP+
k/74malUTSba2G8ucCEYnTYxeZe1zzFM/93qnvJNCRWUXN96Ec9s9BRQwVtjkqMfx85URr1FAWqn
EQVJ+0MPFoh3TP3chpI4S2xENs1UL1utlGOhrUlZc1xciq6DJvWMoOUz30tnCil4O2QMK4mpV8/R
a9tiqU9+aFDChZdpFmcxz26jf9Pe+OCliWgdr3OgE77qfaZ8W/ULSAWaxFJFLeBjxTuac633jJWA
L9wmNe4s33ga5UoQ24WpfTObv54cz1kZEcI2TWRrG6ku4c1CqLcgoKymqCuYNajIfE4na1oYOqSO
fBQ7WtCz9q/mb7A/uukUe5a2/w8iUIOYfqnc7arQpt676A84cDJAkVXSS6xmRIgvPjEtzSmdyWEd
r49TfBaP16xwSj1xKh1BIUy91XW6sc28NmtBiU9bcsT9oK09ynF8t0ia59Vy//0xaT2bKs65wjm+
WedVit/ifL2TttfVy4O6Eftw43P0HPhksEo2Ejpi/BdZwMqYB4iZUhrrQU6JCBr7gkl3tz+3jhr7
bZWsJRlxVRQZMlYe8UZbRFLLhvHSz05W/LBM+/VlnRDf2JcfueTJFKlhkBOh757Tq0KScUi5dWqu
ZV2StieHZwCkYwX0BQbw+/npwzP0i5/XwCfZvRECI2YpqDdUFBdieh7swYyUIS4bIDsUfDOuHJ5V
MtGI9iJ+nWyoLSS1cevEMBwjJOk9pOXg1wD3Gr5JDXp4JnWLkq3FgKHh9B9GxgIla+p4hpCPfEp8
apHpb+g+U6vHDX6Kvc/l2+7E27rTIAQytuJ4Ag0gKGqDoPlJfa39lSL8dg2J/mSvFYiyFjtQ+pTL
3gcPnu5CMl2zUw/4yEeRGnqo51q4ddO90iTFeN1nAE4/e4wkG4iskpoaGpIIRraqTyKzZeAlEqTs
/R0sro2uX3GeTyETU04NcbyYx/MoQqBHxhGQ4SkBfYYcgbONAy9hT1v2kqCNimqw0kiyaZG5nVgy
DRdOQ0IcZBtwPzFMemUFdooTUJu8PFLZMBUT3AXvU6hShCd4GGKBGctnEKe6f2Y/EYIhpRKYkjli
4AKJfUOBIFzf3b4sp4dfyTXnLyskJ70M+7mstWSGAY2ixyXKGKt/EqPPDmoDxvHAyArFU3A+CmCp
YYBqrfHKCMxVUjD1TSB2igl4u06nuftJJLf0T/F5ol8Bhi8R8ueHHQklzotPlXjZB8aAt33aHzey
xyiBQD7EYwpTe8L0o5JSbG2sEhLLzLE5m2fV2gzA3jvCyddaqT0ozmK3xL4oqRO32+4JvCL89hNs
YgPuBNk2V/WKRSip1JF5aiVbcdK3XLfO+3VtX1kC0G6Coy/zJG6awNE5PpCVMwb14caWZmGziR2Z
D8ocFzghO5B4oIw1yzUm/oSJ8HBat1ufzfRKMar/E3Xiw54va9t09pb7LCj3Jrcrv+ZeO5+sgpJA
r69RODavC2VUnORBpWT91nfoNMMJ0/HUhySAKzW+NQpJ9OYzqKDC0BhLfscINMQ2/V0/gLrlvuVS
UI1zS69akciKhH9arJF+fE5jRsXxo5jDaFZMqaE+L64jGVdR/25KZ0c5zE12SB5ary7kWXr1QPTl
rONCzkerYJdpRRZj3loaCMV4BRIM/KwEdt3Q39SRfmIoCk/FPdvNtsIHuKKxHVNrvMvXMh1HkYbI
Cj5ige/byIqUbZS1sYr0RyJZCDhRU37r2jGCHFyvgQKv3cTW82R4iEXYNCMWOWSf+1bkRisdJmQq
6WcdH06mLCSKzpHalRgDu2Sail7jIkjj2jcW1MZrOL1a3ngDRvQ/a395ZwQtVJxniTrsE6Npihi6
9qwH2jZ7Bqw9WBoaCwsK3TZh/Rj6xbZtGlgGKVMJ8DceZ/Ba2Etmw+obsDqWmtaMticMnBT517Qu
IZ3ns85Ie8sN1La2LBeoKMRN8xlfez0cVGnO32PvbXPqvNbVX6QUnsuX9f325gGox0IHbVypckTk
EhcQ0/HatBJLVOKdMWiKHVFYg9eRWK4r0PkkFsWpopL02NPgIoSdFPHcrzpSEJVZ675AUAmxw7l5
pmEJpYQbHoETlixxHTaSl5/lvcvN0iGmzHJMKMjfO2Rzn2J5MBmxRRFkLIa+6pOfi3M2CBnVsK0g
PYncufaAQ6D3AX8nBg1Kv1Ep+Hu6vT70onlUzuV3yxliQ7CiYXCwRGm3cRMtmwLPzh9iGCcLF00E
gyPvRENLo213b8GfBrTaHKhXlTA5DXB2VtrZRs4Ww484Pn/i2OVeDEDpN4Ajy8nS0RBTgm8NCDYO
tPbVFwZdwS3RAxlytls2yGPbfxBBnvhWJ3vo+/FeHXUreoFqq3/Iu0XVlKK7l9UC6LLDbyVuM3eO
5l1CPkZA+MWJz6nRNbnfTDa1QxxFAA9RcTaQCfgTZ31mkEigX9wmgdIrt5C2Ysh0IDQa9bQ6yxjZ
RyTR1r4W4igxepeRdfO22l8eHch1NwhusABVoaq9kmsUMV8gwHy0wMTCnK3/902ZXWg7yVJB5D4Y
EtX9eLFwXJNiOHx1wMDeQf8SuCd15hdp9of3JToTlLh/j+FlBKcc5rA/jqCAWmNJyF3/DzMf9xHc
edpFfAjrQyIGJ90CrA99dYcNMIpt+bJUQyP3LS/foD+jnSYYdPIxPqd/kHvFx2miLWPCO2xEGwdn
VHBo2l7bSUDFenAM+JVjUvpfe8atSf0xWH15EbGe3gOFrFaOe/Xt4eVjMSob6Hdu4EagpvKfPmMG
aqDG+U8oZIV25a29grXZdRcp11yJqMdHcGLZqP8uUPmpAdJL2yVcLVXawx8jWt6kcGpjutZw5Kaf
jE4kb7LaXTLB3NalVlTSGwnYNUMESlsXGGFnUGe5sXOU6/FqY21Y+ewRru+9qu0sqqGxDkmaQs+8
Y3mibGqU4HzB/nm9iWJZOmAfJqsfKvadkjlJXZxZ2YZgDcU3ztOjllzhXhu/2m59EK+ozBVDHEFG
Rjl4tERK4VKXsLt/AoWR+CNluuyYG8EwjheXGqZISHEY5xHg0obD86UfbxbVZWBW1QWxfi7hNBfZ
jo5cIOkEuh6U/rWjB2iqgwBmejeeCAu8EdWasKQDQicRUDMK3/y6EoZyVzMogHOeDyzQAOOAZQN9
BY3hCncTG3tLuJeVECZttGD/OVXd9fSnPiBUIExN/0RJGhhTgldztO5ggxVZxyVAKCEYytf1zirb
aU2ETRM0jRXLgiOowIbcxchwRvDAhB7JWg0N0ufKrTzy40YVuSxyF2WNLex+Dig1sxkhqbgs6ZCq
xBXVPai0q9qnGSiRtzs+uERpx1BCZJX74Blh+TpXzfwwYtahC7hTcn2mBSPbegt9fz+TX5JgtR/G
qgm1d0v7VuHlvBQnBn6zpsATmx57VqWVg2t1Z4n/PnjCH3XcboY9bqGvm3rGWmETv/FDYUHgIU/k
2T/aSuPB8qtcRgs7rwJBWjZ00gMMSj2C40Agef9zbyCqzsOZDUQv9ZZ0usolBZ4xXYsnoxF2RCi8
g3glr5hcUeVl7I4+acvZ7W2vs2yQ0Odg9VrBIOCoBwVGqZmK9dOoiiX84bg8soosJOnVTFYuWJP3
lLtws3pmmIue2+iv6HYQiiUH43T9FE3n0bzPT14/5UkQNaAS7NQvgK3GA23hX98bmFoPNuDEfYMb
RAvuP+FU4zC828gMY6lHyl8OvlO2nxdv1D5P28qLRKSOk10g3Ky40CoCFaXEum5EtXN/WhSCk/JA
88EgxnWG9SOgrI4FxvmfYaToXUGY3EEEx0q7pA+k3ueYXbym42DpQ8B0fd0ETGRwO2oocAlEwDjt
9DN+6LbVvcSWw1GlYBKM8PwUmeDGhfjxcxMnKC5YNscLQsmEaT6vvWcFBUig9QnpPLtxk60pVh7N
2FB8ghbAxbGZgY5Q7VNc1/JdmnUCqDzXW54kucQcxtWx/BU7NDjA3Sa5ZrSsVJ5dd8gZbqW/5+PD
F0a+6GEhNWW9UZGnIqkq9MwwPkspbDu8kfbh50QW3fzggE8p+uiVF9Xit7KPkieCdUuWXkp8oQio
ygHNDuO4JwXJAXmNoBaY0wmHy33YgVB/UC+Rzdv8Ie/jrrRQWncFktsI/i8t+zt0gJdpvzbz0UYg
Sp9fk6yWp+WE7u8Q+kSE+XVfT4clSijxDOkltEl/7xd6QDF8FwTFnLpELdiSbZPV/vkPadalw5jJ
soBuMsOqDMo2/d+anx0bnrjtd0P8t3Mx3vOdhg6qOuIcSgTAO1N0hDxeB8q5ZdIP49J3sDnK4Hmo
Dya7Gv6o2cj8sPWhACK1ClqPhMKR/j45pAkP8GvJc+2K4i5juDOzODvYXs9cOvcX1DDFGs0ezJSh
7XQXyOvOaFQaDWJNbfX8HrO517ZEW1qAQ7mVvYaypzZvsdL1uTA3TOz2y0rGzaG5qfVKB5vls48D
a/i1c7YzhGdv+xS0nUPvzCydZAiebt9+iIpjvq9KbAX/2mz4zr+V0ThVqdRVjn5LDkU4fVgcwR2j
nlmqqz1YhHwe9p7xJc2S9eQLY9JMqo6hsh5TroawAqj5ajy2J/iYCbYmPzainhoxMUn3yfuS0TwO
clIDZtVNRFmPhIVZuLf9NKqIIL0EHQeHASXm2kGzJbAvAd6hZaeW8hGLOEcMqHU2yEi7TLvf83EU
UM9DRE1lCnpQ4gpcMm7DJJQ8P78qQ6JieJ80AS1z0Jk6XIwdr4Ka6fhAYP1vsXj9U0pZZnVYwxxc
c9LRU7m7icPU4ln/MXduAZ4WgZXeo6Jno2iOc1v1UuN+E5kmqRvfCNxhLWHN9zPfeco27E/32ato
im/cviCiQerKD+PWSGsEl0fR1h6gM8YRVOOBFEwzeadOXLWaHrdijFM63PSg1nHGrCcUyYVqDmED
jbb4rVw80AsQsRqXnHVhWvPR2fw9fdSLrtfGOdDSTBM6RpGJBi+wiWgBsyZyp7gD+s/93SXR5zfQ
rZELhUliMaNXm750ZQ3cDGHjIHJTyqZnPFC/HXlOl3SAmd0PJG0VZfUz52VoCNCIZsRBIcT7QuZm
pb/nnfVL49jThXgoip3rvLLkvOI+vmcTm2cMpNeudy/5BdrahiGFK1UvbC3WdHUG+Q6xpqGMx68n
LhgsqpWkkbXgebJ40baRrIkQOB9HqtuoKDHi8ckyTE3gpE2SDZbqXrSJWF/d/Ds72MGWGpd4k97c
dxiByTMQ2drBODjj4zbftuQX6m0rkAdfkcci1H8bNHF+eTspBcVZen4POVVwnse2NtADM/1TeSyG
aBXy+GY0ZdB9RI8KTtGpR7Xt8xf814xIPepdFBBYHh18+d/441sWAWtK4y1U+h2MgmdsKT8Fbkma
ileStH18qck6MDtSZdTagCXcywMZyJZZ1FNUwXiARSLBs/ALEtYIfkHPgzvT9lZDcjbaanasho9r
iDEsA7bjHdaHfEug3irHmkDFy+gLvGtDcDJ6kONFq0p8T0H6O9raco6MaHlRsABmGGLPKBKA/G2B
xzqh3trRe1VWT8fvmqQMTybV/QD/FXOSd15QNEQIb7Vp2ohzSHpGcULMbTQI6r2nGtmSLsbwzrjD
DdqhE5tg+EsEUTvM4kA8x1/dhU+kBzO+P5BW2dtLbe17obSoLEXw9XpGJelowsql7Mb1EoNuxZ6G
vrq5p16XB6iaKSORdRT8eIPmelCRwlZXGx3YSMOe8ZGYeYN76n8EqO1p5/B3ob0T2E1lR9Xir9jM
XYOR4SXXPLSeQHZsNv3FJ1bVa8vyj712wuxPRifYFjCmuhEuKc6fAbwiGSyrvL8cemPt2VLm9G3D
Sth+IoNdfcoqJ784XKJ8H7gyVTPoHvnlN4kgu3vD+y2GuwYZR8fAWF//uFoU8sUyxu+9tt5I7qmF
q2WSdieUbXRNGy0AFqaJ/egFOqE/bTbM/FoI9KH+ABCmBv3Bs5KddyGCGHqrxYUSDeqowlAQJScx
UD7+1Vmv/kpkLzmyqUd5uI6E0DqqKKSs28kgxRYlI22T0a//uK0nkRB/N+uCK+YxPj5ghcE177WV
GUEM6tVTvgFSksWj4srnSj8YOeg02aKo9E96BV///uxzEiqhdzT1hrGc70e3GmAeGJnoXXY9j9me
7Kf/Bs5zp9oFcIyf305ekgMHvq24jc3wNqeLodJiEE0QtFU0Gatxy7n+5Xu0fH8god7BqdcsGsxs
M7tHhkrw/J7O6/FhOQ1XQ7CcW+bb8RxeAj+xD3+OojcjKhwBc0E1NQTINvUOGzzSdjOkj7BOzED7
L2DGYEra3QdOAuUR4ykRvFyjgcM32w7dDAosd+oGZ7rhU48jKx7YvLBIR/CQCMZRkQQ7RHrdFAqC
ZWGO/lLbEBEMbMJC4b7WXWCLZClQkJQkvKls8nuI1PMfV+Qpt/mgO/9d+mATtfckViYSPQXiNBxc
1Y9I3CUhcjGvGgfWNNJdR/p/oHqbcGUgopEi52HcQD+D+B5MyqYpOjLmpreuuq6o4GJmYQSy1Tq3
ozGry7tdGHG2RsSnPlFVaQuRKJ+capyyRfdtosAQ9ZVnlHZ2yylSg7hD6Tjvp5HE0m1Lrk9dvdgP
zRF5QXMHWsoxrANyj/hCE5lU2yCOBoB9s421phcihcsQSdxAll+F1DiR3PPE74SbJa9rm+T5Dz9y
Bnr6YU5Fq93UZsXnw/ixJjVssBbBT1+yZZxl9u0ph1tgio0C4zwL2qcNDo+D0QSqEYqGr/cTwpWM
MN7eFET961DzCDwsNrBt5GGf8gyrknkT+dFAmEfASusqFsqBD0DPWisFNsBKXZKM+hIG8mcgwzgC
bNQCzesg3+DKls94DINV7lNq19T/jrcdmr3qIRJa7F29bLcN6Mz3C5U9L1BNFa7cwVvzu96dcOM7
1A6rYhsZVP/p21QgQ4NnwcuU1rihCPGFMxxGwmynlx+o6FFXIKATiEdj874dSGaZQ6xKjklF/8E6
nPXuU4jLuXhVBfWnYM3+UXupZIajxj1dVFViW8aJ+/Zyns6vFLzcZGR7cbaIjNe+1s9/qagjEbJX
rqu9nvzxZUfBI+TkwFsVJUJxsAc7y6cFciyIqmWaKgpiLvp5FoaCNZitUn41VI9FrIpZyh/MQ3D9
X9mi2rO/PgAoCg0DHLFWNDYA3WkK4LVtNjaBbZXSDKvlNW1zfxpgg5kQlAx6LS0HPxZZ0pd4MKCr
CQYszc40t81qWM4o/5uiT5ugPkUJqekrEdyf7PhsMqVurLQNI1tnDUd3efXachJIFVikD4Yv01bt
LtTQALELQQfRRX6F5c3Nuz51rsnvz5CGuCBkyldSXFL2euv2QpLttDiHbygZzZhGILXv8Tm2/zBn
NnRA4x68Bgvq59Vbu9IeBXWWWMSS8SFPqM8uPK0mR2mYiiqT3DqzU8HTO2frLdu+BAYO5TJSg0vA
EG7auqmUPiAIyGdhQR8aOiygGbpZo0Jg5HS7ZNXeGBhW8pZ88PN/sJK+OrhMeOAkujVovv6dlzWC
wzyyYhkZM47czXMKssEHHzXbvJOnrv/oKIgEIm0HACyOKcd3frWrVRfVulij00ZuyBWT3FC371Xx
Lr54pHU/bciZ9PdlLRQCkpioKpJS5ScLnPpTzJikdLsbDwew3UhoTWvU3hAX/YQUhB3JaA8COBcx
RDmqCgl4/NStaXOoWRA6kbzsxV3NtHU/Xmkr0EAfEN14++xZjdSrq3Rd85HmRa5crdWye9s3cEWn
bngz76Ja6UGkZ5tk0kMC3vmW6kYShFlve8iHoAVL0GGlAOzVIdWAvKMQVBUDjn/5l10sTCfjoGbL
dVj2NLy172LQfIBHDJu8j/eYS789IMsvlgmuoO9xWSL5TCowCOEzIT43ycqq0bdu8v4ja0LTcEid
JOunb+0V66lPw61hy45nSJba2va95+8Csjo4r91Tc391ztx+/9wXggIvZErigutwvxJHm7SRa8mi
1s65ahsNhieEoN2b9jb4vc6GQryply1CNiuC1CIAJMpylfVqjUyRE8eh58FUnKGu2eyZK2H4vvMh
z92A0QF3Hb8IgvQCla/4y6lxupksQEwzHQSi9FzECoAOxYTnm4xlDw6Od3lrYTqK6yMQjncWVk5d
T/7jQ3o7pwhwiMr0T3QQ8y23cG56BFHxFOxzML2lIbMcltAsNZade2WKGsz/HJb/0drIOQzPGDZq
XiD3QAyxR7gJOPeIlCGmxB3NuQ8B6xJjTpDlmYp8qVMbsv8NcsWEqTuzLqHMDF4hWlTNKWJDw32j
zWwAIRv062otHckPtCo4uFG4Ia2aWB7Ads/TvUHKZcO6Q5e5PUdlkbkyni6FcDHvXf3QTUCiFOZx
rpGhh062mJfUH8Jus25hbLi/aL1VuH9LQzaLmhINN+d6JyejtmJtmTipOJTFxuuil5rX1VWL1uds
X35n4jRcyP424GDqhOvtpbAbNkyh26V437jXD8AEHxTUlyq6Qsj+fZ+YbUeZDAdvxH2q9PPEsodC
d6Y2VdpLZ/rhz0xjuBcgNTC4L/ZLG/4Fl51gZJp15Cs/acElGk02UXf3Fhy33uOexz4kBsOtfDK8
fMXgyOGVVgvlDGaUOxqYkamwsdWURZ9xrJCL/dMcPApTx1WPqYZoB21V06i2sPN8U/iOobAwNJ8/
vYtSC9DQ/EQOg1XQ4SZWJtmyNRwF3ZrIT7I6PCIG1UuyqGYP1YquCZvHStAa3GXA1ykXKLw7ZkIn
auU144VWZaLU7wcESGpWhdCTFmv1b995hgsEv5fCjdvJXvfifUqnLI98lcsKfuj6SPoqGG8OrwiZ
sdeQepCTlG9NYPdq8iNnbXW9tGaKOjsCudTfNl7Ovx3dp1TMCJhL9sGI2xcHSjoNndgWnZW3W4rU
XbT42sihyvQYEIXw0VynxfGAiWsfpBqb3xha3xyERD8ej7CNfZfg78sVk++jtkZSPpzNCmFYVSQc
mL0tOG/BOFeaRDnQMA8SUy+N3udmQAEBNrBcv52Udxe9r+BBbTK/7icxQbbyPTm69IjSRxNQ4quk
dGzHQN3dlhylaNHf0oimR+7HmIK3glvjtAaj3rGhiMh9XlxAuL6tk3llpb61/MqGgW+LaLdUwEkT
TCyTlwfd9XGKv09e4DcZxHHTo4P63SZx7BWvcLHxf7EZwzXUV1MrZAR1nvWqWyz5kRUpQ3SP+2Nq
ioNi1AeORW7TZGsxPJ/j6f4TSoDseGmgsn5WQqJRK3DZs0SYGOJrBgOVUSHCXTj0NOi+FK9YxCuj
G/uoa+VD6IqioDEaHtzlWL2mOX7+Hsy/jzvXWL7rTHZXxNtB1iydKyr+CBuA9cvPmnP54l5bGeRz
062eT9R7XEbatJ2vZvOrDYvPxLY4FxEi8QUuBrAIj2MevfYStLGpLSZKp398+C7Q8oejO0F8fFBT
DJhOiJ6c++BpFbfSW6CjOeqRTYj7o0t9jvEiffwrF/CQZ2TLls5lOwd3y48cUg7ImdECUmDZG7Uq
gmrFDDsDI0chZCIbzkGIfk04Yz/+b3bvKxMiORPcmbKkNOyBq8xBw5G88Ql945gjMCiAyGObzTop
9xwhXsg86NCEFOqsVcIpn7YPbcdbZYEfWkOjZWUOosxE15ur9SiZ9OKoTXVC9/EOb1dfOWccte0v
zV9RskEJPA4608o9Krkkmy9j12BV6IjqNpk1tql0GN+kPyEDKZP4F3VAD1Yj3wgTrzCpWQReBROZ
pynA1FjK5nwDBb5qXqmP8MdrE+hX421IKMUReezTmHm78l9z789JvoPPZsVyBa/C1ZyO+c62So3x
h8LaPeLU5SvcwgsLqkqen1tWJGAV/s76SA8YbPVxhK4k/JoMiqJzWwk+EMnDnK4zJkrddyKG8xqd
/99G4sb7Fky7+KMFLJH89F4ciWLgx9zBn5nB4C2hddVBdt3fmkqrUWSpxefTheG6kbgevpe04Ail
jdrC2aYllbdHfxEfZ+CQ0O1jg0xRjTtxtItHRqiXJBnceZVk1BV0IDhxUNYZ4dDKBHMwnRwH0QfC
R+EdSPGEOvoPzoXHwiiJ7JGJMJPLvQpR6ZDHJp0WvL/jJrOB81V7N2lvkZ/6OP/7i3XaieD8TQ3/
NECTkqHn5xzWXQS10Z9/UHP8ki8NgxpSQ7rVy8UstAw/OGqP2/GTQf1Awdg2T8XK2hH7baYpo/hE
6lSK5iPws/rAfjK3z34SlW83vMbytMJnKeWypVrTp3/PFatVpD11kVz7/4t9BSgY5RoL89b36iJJ
axT59D9W4VNxI5ZJ9a6CO//eowlq8bSlTL280dTEXEho7vJT6Z8=
`protect end_protected
