-- (C) 2001-2016 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
LKlITFDlw1rfQMsm+oYU5yaS/wjYKUhl9njtpQbH48jMz6IG5VdxF+joBSpKTcrT3Vp/DjTSO223
bbNx7gEc3Aw7C/t6+EHxF4fAyVIU/GW/NrHg/dQRD9SoyerFe4YP+YrLLCpa9yFWWhwOOvnp6Ldb
PomAc1o7mMfeypnt/LVIaydu50J8IelfIH3NbdMYorCUt7vdrHvl7A+QHtBpXlDFKgjdG8I0j/hU
VtUD/XL7XiW6cCECcWZz1kxs6Kb/adlCZfvfCEE4/HZ6z0K68NEViC3q981nfRWwBiYxBhnC6tHC
V5zFyYPopYhxff/VdveOfhW06AW80LFa4WiBmw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 10144)
`protect data_block
5QgFHAxZqy5Ll4V2GYFsYgKZyTH2E4MgIpu3vfDHJtB6wXUeRqUhW9R5dHwgQ0tdNMN0LPzNyM6Z
FsG8Imc1lWc+V5j05YD+Sul8oXFlvUD9S0NmiTMciUSKQszVe+9bOlNe4AXbFe/EUn2s+8HFvyCz
f5Yg6oPX95bd1uUUwpepot7Wh5OgNOJI6IdWwkfGIfSsr/eB6baxPpkLodaf2y5qgO4hJE1eUFuI
AmZNqcZ6iEvPFD3qLU1f7lCokeudRaX8+SUloLmyvLRexXuyZYrjOnU1SHg+CXMUza0r83sbTCOL
sTaiYVmDS0nwqfmCOAMHtHX08C3XGuG2oqvpRfz1mmMq7U3zoVk44kLtb0+9WcxptUMahoAU1SgN
I9OPFudQl1GxiyCOyZ20cM6fwlpKHcOKubkw6pA8hmv+Huv4zy1wpYpmUdiUJzv56L2FaZ6R1KK6
8KePAVP34vazhYeBhf/CfB1u6/pTVsR0Vwp6T81hS12C5c3//1RXV+tQi5RhAWSDFzUCr2fjoVQ5
h5uy9ckSp2oXMwlpoatbZJHQSa9wIjp+zPqrg6krVihKtJPJAGjdl8BkjEIR3LqyrXb96VIhg5Tx
oFF69u856qnB63oy/4yJQgNPY4VAh+/dsKSB6U6X/BTgic53H4FZELktTp9zgWW9zJRhEkBi59WK
Cme+yEkyquRD0wmCugoY4z+9efRsrdgoLE4zpAw1p6hyat2hXT9iqozT9iAouWIkOYzoHxEKRxEG
I4QaZw2xAaAnLP73msBKJviB1LJuyDAO3GBP+vVwRkX2rU5vMMTMAI08JgxfKGApBqerAW2+HNxb
c1AvUhVGWgjXvGI2GIbJ5rbwYdXT+ULr51u0qKHNCa69+O4ry3G03LboNaUYTaBzxEenrxk2xMwb
qmtAw95bpfpFp5X04tAGsHY8TP5uqfTBi+BF79Bt1mUWVTxG5S3kgEIOhQGbfsvt7a4L4vRvWqgN
drX8i2y2o+NOZEMAuCtjQghgHTdkFOPX002vWEB2G7/r4LVRK+94A48YUpc821NgShFo756nKsM9
7T6zgrt3J7Bf51OROiON1QbX/0XoYJF06c+x2BJiM5+xkJw/k8Dk5WZ2B0VniF8d78QJCrBKi6cD
OqI/RdqbC/+8qYhCCcc5kNI6pV/a9r+eqD9FWfxVe94C+Bzs3CIxWB0v7OO0OeEASBGhBt+/9vww
8hOqVBJTfyi5BMLPU5DXJIrzttDLWEtgwo22NeEhLpj2cDz/iwVgumaWoAfzri4erapgeNw+XS8z
vTpxYulT6GvEHA4cD0XCjwBuMm0c2eH9/88h+8KJ6vwWfMo+XLbvAPYLdtgkyF4VfrS7DRA5y3U2
SiT7dcKg+5HX9PVmH771uShT2fLW6YEH3r0JLYqIeVPHp6W4k2NB7BRulWU4qovvRfZCIREonhi5
QRP1exgLoYXfutnxq8DdrcObfSRP8feUOcbXLX15DWxRCknzgB6JIvfu8aiAvPVC3JfMWVb+Gpbt
kHe++UEC2A5f2bkj5ntiVrMI9BaR2nyZm1mLaQWWWfDMrZQSk4hIATUQYlDSkKqeasO91UQ+xuuy
z730AFnGQ5ox7XMBj75et7bBDu1mwXeABH7XKfOY69DaCYKkSuE1sDDJ9IcemxxvgwxmDehWa76F
QrIq0P1MegFP+oqomRU9+KRnUMMwc2glYLN39zwdp3G0VgLRexHlYrhQGbSlOhQwdpEKaCkEpHpF
eMz+Izz7urcmIDVt7cekg2dh+xr2ytHZ4OMX3TBegyonaysAloZbKlmuAkpjeW2hy6hm9l/PRfeo
il8519V2m+Pr7NzJKMJwp2VjeoSbagTy9cYtX7dEVh9GKTfdYSsicy5KtBCol7+WUH7/6VyeY3r5
TUPuKyCLNnhgc6dN4DP0BcAEO+WaFOdKtob0Twb93MmJ0yp/agtBYKIy3ved3Fr+Dw78lqDbWNgj
lpS6vZNgAvjjnaU6lO/JCfRCCiEcH0XhY7f9IXjeNaagV0JHP3zMVbDc6XgKHzf4AtG0F4mJbajs
Nx/yCt0oaLl4Mz/KApq3AF11S9jt4zqBoQMKxS8l4QAVdNyBnBhUhdueIaYcX5wJaGfenYE07I0w
ubR5MoNQZc1TeR3AL9rS/eINPplbLbRpM1SxYV9Al5KqRWPC8zUxPxUXTv5j8DkRTLREnoACwwk3
YaE4Q4XQgWRaXj1W6qC6BNw31SczQ7FaRqQvs2rYQiwk8pXI5a9Z6sAZP0LXUzOD3UtFLHr/PrkO
jjo7Z7b/jK7+nVyltEI+I+Wavvedm/+4mMUvXj/lvmr8hR6yr4sXDRyLMg2+ErNZdL1fJbiVX/cb
tKTKS+C/p+TEfCBbTU/ru98kwDdO7v363e0SiYqXJFXtv1RBWPWj9xRsy6LsckW+wmW14Zll4c76
spr6fTv1rS2qsbghAzdx3pxXc1mZWk/6yi43h2KvBQ4IfyCXP3d/sZziokckpuQBM6FAPOtVjeam
OaDapKz6ZP9FUE5IeNcOMoObJO4QLJnptafr0KfUDNjc+OUrWhvoe0ffmWj2cqdRM48szVSoyk4W
J3c2GvQKmN9nJ30ONF1qHhVj6mdKt662ASrCZcYdhWWtAkqNC5Cc1THPNRjqbTVRnLp+gvx9O5w0
77k6RKdYdz3MAy2rlf7Igxmya3VZf38R4xf3PmHcjv1nJ4W7Y/uKKfAq3oyBO0gzuDS8o9V5K8xV
aJVBEcVWBgj18Hwhr8HcFi9x/aSeYWOLXbs2dJ+yM8VaG4vlXcLVrmVTk+YtRuGI5WFSdgAro4Ub
3L4wSj1oi1at0aiO8uydhUtUYaQKP2f9fmf+X03VCVjzxN/+6fxtgfpehO7TXZA47iXvHRmRYsG/
pwP6y1b5zb9HrgWTfsMVqx3CGUKVw/7xBDSEzzy0GjcvQ2BVkSoE3CCS4Z1YeGN6NNJnXEdIvMtu
srOSmnak5tZmrLQku5TyVYNbk9zzZBmidzHpgx8gfdRoyqoXFxrlTA8FQSluB2LInqmZaTmkJ9kk
3FPVm/99a7i/DgNETbGzfGTEBIsWVKWi7scCzvpl4n5veasxsRJZGkrGrd9a78yF3wQlvNIbdQMH
MY4BiqyuvcPbi39ayblZCiUYx6WD/8kGkwXab5UkE1SuJUoQuld8P0QgiIKejPfm1JbaFYHWZ9sN
tdZgGH62CD3BIZycGHpypayzmvB59ylFIaAYxAKh0QTmBnSRQ192OtLDE1y0uldJ82P5EJMacwGE
o1rZYRBJJCsraSARDSrCj+qONDOS3cRwYtYAN5a70yiiImQHi9PJCCL2V7tLIROmjCEp1DYrQMAd
hI7ygmO2ON3e7Z3sd9zdKxeGHrg/JrmhZTeO0jA9BOf1Bpb0rtdSQYa6kWhk0NiQLwGXuOIG2xx0
wz2Nkn9YU1LoiV5SOsxa10U31plWVKfpJRCaIrU2kh3tsYpXF+nvcO5UWjo40C2pw6lXRraZfCZP
QcbOLk3kh8hGbn1lgjrNQs/lMSpa5NpfRpPJ/kthD7HLIto8nvojnsnqV4kdljlY3yUDnuq2Kv1v
BGSr966tX0DpG7K81Xg7zXh9FDK4Fxca7kNHs0HAzRWp5BY+vZ8HHhhlTkTQu8fEUPnepcXLn1ba
b2gauP6XZddqnpbTn6PbH+Ow89B/8VNU8yWbyfu/GiVTlaWlaQDOVBa2QrJ9nKMzv1Cr2RdWcMhz
YCflpkYPS4LJpb3L0Qw8D4IippCyo46Do+eMm8kSdCTw/lIcX8YwdjELQfgYdCpMKEAXBPPf+Bhe
MIuh43Husa5P4jlYBTc5Xrb/VUK4xmRXwx9OS+PoncBWW/4OBmskKPRsRw8XpQQNEl/CoEJUi7Rz
Aqe8VdgzHFSb8Kf49TU/1UJPauMS24gFkuCpGKz1LJi6t7S1uSW95S6GXcf+BJdFk2AoXhlUVpVF
b1JfwfOWFKRdj+AYsOP35vWSS57DhIJRgRdrUYC+Cg5/f2JhbD73ChSJTasTXc3qCF/8ee1JwTKL
NfjodlFQype12BHfSxOVXH6ugoBSdpoR0WVXkBbWs9HbsKo7tuNjja5qnCKdnXvvg8HTsJRepeGA
5IvJIwN3TrUFy4A+0N0uA+9j2+VZRvDTdCrOcwmmN0isPs13KvD7QY+JC408Oaiiw1ltTELhBSbV
sP3hkc+UwYNsjy2je42OhLLomYrLhnr9lwrTHcBrujIiAFp5kD2UnJYOpuszX14RHx6yNYbzRuvK
qeRMUy9fA2St1P2J/CT+xiaybDJGAzMGcHGScTvj4nGoTM6TfkA67T3W4812Zfzv8dcAADgjdhwJ
gg153SLrhrzHh8ahswN6vAtmJxDGv+2f/UGsGUC2AAdVWtSQDlrPxesokPbEuuobiztn4XOIcY7n
YrtJKeJTK/EHnVBEq8vABjv05VA/8XZfu/WxgXE8BxNOWDjg5zcEU007Ax2L+V/43gI5gkKrQkHq
pA9yqJ2+zi2u42+RNgYjggx5S0U17TZMDJy+BwysIEjo1gKKDbBxsFpGhyMOJzzjXf4hYSRba7pA
SG09p3QsXVqO3ud8jFq1i+5Lia53rB1DdGgOhFeLGCtirAggjB0eyK3JO/ACiPOHYxjo76SI5iJJ
TGs1kefZooiaydejihtWsiP3xMpCsWkd/1qliEX+HPVIZbhDcd22AZwIw71oroSmS5NXY8kISPW6
frs/BcDD2QQceP/RXmTtvArP96BkYqF2uJRbDVkkEiYnwPRDLXgmi7zO7IHm3QFWLsPF1G5LGg6i
ebyhJDPNpUpul5ErPsgMoc/GRrCOshkF9pd9+juu/678QVl9IW+xe6zD7Jm573ePPmj7Cie2gEuJ
D1ceUDvPjbmSlu9nc12GtzKx0BEqyjLlnO0w80++sviXWAKEazIJVuWP9XSD19R4Xg+n/LZymaqs
V0RO0KmhPXEL3aTxHh8I2ZWoIDHSZkq5OwSw9TXIYO2xfq+HtLZ3FHH8Qi9RvgWLMPucJCZGMl/L
YswxKJq295KmjFlx7iv15McSAIG6aanzqtjf8F3HNOKz5kju5MeigFfC0gplko3+uEOxgj12VK6e
uWCfisa2xVnQJUz2Yi13hPw3TACj3quxQG8GCa1RGGmU8XXtykVFCNYfe+Pudm50JtwPVIW2+fyH
u87S1M+vGqmuvulHpUDdgLLpqbGP9Esiuy9PyOCXWhsGQzhEYQSFO1ayQU021bDiSvgQBx4uL/Gb
/jailzeJyqRILl0TOWBvQpp5Di/4FKm6n2Pzf92reZeZ/BX4xW958ZWk7ei/f3pMT+ylwPpiYOEA
ab4hjcgZaCKfxbNps+5eV51E7xJI3qYRHuQElnXp42yKi4PVHVtWjBaz59fBPKOs9JmKPg7hoUYD
A7C4inHVf9e5D0hS6Hlm/Wg4/FI6kALgWpC+ZQjFsr5EYRSBhrLEB9gux2j/os26Fi8QaGmq2zIh
fmWihkvc0f0wT7SzaKcjPJStpHIAlr9c5rpalv9Pzak7Eu0AvHGcZe6RsiR55RHZ94WLw0+CFGg1
KwHRrvBBoe+Yse71xFfWJUlJbnmGJ1aZN72GyIXv/tqfStDjvLUksVvP68Q1fUQNP4uBOYSH3Pea
JX5UwrDJ3nuWhMcXtDBVdV1+gQ0LAafQDJwtf/h+4GDU4j2ucNszNdKRfyZeO8zdZFV798PyqWjN
vPExEa9ruAJeE2+4yKatjccv2MxwTGpTEw/nTB5+FIkEOQEIKMdnVUkg9U3rtKIAjnaLoLqcBQcj
kEeFTHyselThbaPjQjgA4gI1ZxxdB9DPMLBT8d9NY9q3ixqVryLVhfXuYO63TafRPBq9Wyk5izUo
YuX/2vMS5XonZ9iumw5Ey3kZT2BG8xTM6HVjQdXJzTObM4wTY1Zsd63qC5MKjyCMS2/UHVjMygcU
aSnIrnhsR+hGRSvjUBeatIfNxvWR6iDQlkTwUtEphXXMMFrz+PlLzxqJci//flKjbCGxeD2Yl62I
nx18ytM0VsCOs8Ab+2jKikKcQXHI82IDc1ivb5uge+wZk5BaRO7jpQrxAbRKnO1KKOF8eQ1yOUBt
iaAnawaoJtbZEwMGpYpaiMufZ45HW1WJ1aKv+ow8ZkfQjc1Ursjgkz0C3WcC0frdk7ue2E1ipfRW
iFUpf9Apwcc+WNr0LYxb/pXfA0Rfyp/Dil9taCZmmjPsC8wjfOwt7zNAdgrZYmra+qvlRqm+l9tc
WJNRE8tnnKUlKwPOCCOLN64kcDAu2a0E9BIpFHg1fGKNBc3liDWsG2vXLo2tsvcPQZR9RMXBnwxL
5pSPIP/1MEtiy7oRRoQhSp6lDKFK1SgvQZ176x2f/lqP1QUykYaUuGx9cxFWIEBiMp6Urmgkkhqe
EqLYmnC0x7+ApizTIWYnXyyfiIDAe+bgPFejn3k0TggXZBLKnBA//UTRR/MmEnx/pIAbogtOndaG
EOkkUSugcOnGn/hXu/ykawQBJUO2VWRhDKa7VJarXcyRMx5BI0n9UMmane8AI+TUVAnvZ8lqAgsV
6zm0L8Icgp6LanJtZ1wBJHFgY7K+ZY6kO9/Q+tgIiMlKaIq+FFsm/I9Bj5Uh1NG+6HJT5TCkcxc5
kkOjCmvtM5mv4n5+HAt37RKkC+w2a7KvL3/5HetP/7DtNqeEUxkheMLOgjak+iyAm8ZEbpICaNOd
CWo1S9wCb9qeQ/LTpkGK684k7wdGhITvuRnR+SnMDIglxGRIijQcyzrWi6uU1zhyy5ktFK8ADwko
GgKyTaEVDiR0ijipK78/rDrsCEle/tzGyJScK27YsjlTMeeI6eCsD76aXiM4Ju/ObnfRuWAqWCD0
cyb1Oo7mh0puhzggsdDsy9St4rO4gFxowzgr5Da0iNpR0bzOUJ3dhHihPwOsOw32FyFYH+4xcqCX
s/x38F5Fc1qwpXnYha19+M/m20URz7UiH/20bLkzlm1/1+rxVU8jIxT6i0MQ+Nn79mcz7gZiaRVb
IZ1kA8DErkNJi8qTEY8lFez00IUi+X2HVhXDdj/jlD68rVl9NgNmeitIMmUCdePxNU+TmbipCaoo
DEabMlhpgM2ClUf7Oo5lpeG0eSRkd9/UYWSXdCqaQoLVsHPXgPNqJYY8HTsiygrdTH55TfsosbZO
8RX1dnkUBS+JhxEeKWO1jlnutw51msgOp+taPeBO0lAmmHqCoruvmHrY0eb4Od1a7M6LcGIvwPab
Y5cedesRZJ6sm3J1Rn4gU7w+3VupCEnPmxOA1OxH6Wlo0cSZXiHm/vS4UMnAw9PUWYygx6w2VENH
sOxt2Lk2cL1IA1J60MIeEfKg7rdFAjdAmJgW7zAnuboneOWtoAm+Y/twSg/cSv+7Wycl4yQmM/ng
buibQuJo6I1kTgZRiBFPVfY7NtivdX8j7fYVknIf0QDeqCnGNA50Ddaq+tg3K/oAs10EreLTVgI7
UHi+4fyyTrWo0sr2mnp/Z+/5p4ITN2TUVMj1tkqzuwvao37XyWMzf4a99z4465u/s3twbEu16Ysk
Th+SXnGTmlKrafM6+Eqffs3lr87LCFfzzXqy/aVCXP5mSlicP3T7zsMwEEBy65fSFa+rOW6f9xlB
b5Xi/83nCtQEPkvNj8vO4jCOqsvlb6k+/vDQA24sNJmHX5OHpWnr32ddB8Vxz8x0KycAmLkS97pg
sQoAMW71Wl3oc6FJHhirRSR7e2LS888kit6j87HC0meaZwijjqzJNSreR8o43nSGcJ7AKFjAZNiG
AR8U+eXm99q2t9jfPpev50nAfL1FMmXVjGPkzZDtqFB+EJ629HyfStMMi5ZQGEUxfwLw6fniNAzu
+3iEp6OfLq9XrclMHTyB6ufmUOV5/ggEKZU0xRmQghmrtcWBl4AyxiZbHCxe37UVsCTMrcVUDr/E
9prPNSmbmMbda7RP757uqfsZMv+274iSPDRcqRqmAreSGjQUXi7z6Hw0P2VcOC0sja3jNRNG3/WJ
HHHMp9VXTYVcaN5AE83abGhDkxTW6ApcDineQB3p2t4/zpiRNDj/zTnZ9Llwwhuh+4EyN+9ExILc
Khft5e+OQCyQb5yVLthpy0hvLOOUThWx0ExF/w+iNim+R1nWO9WKYvrxAfrxi88NNvIrnjUx6ACx
Wt5H3nHdg7QCNCIeUCEPKpon6w3aB4pJ5MuybgLjdzwZvSQxSV8bQncot4UvbPwqnbrKbw9/8fzi
at7LCdCpsF/sJQopscpHJElEMtPDZnGtNQgOpsg1vNBdZM2A+obfKKhPYbVNkzaWPoXCihjMHlBe
0uKPxkOPUVGxcrRsIjjLDHsC92thevpvQd69Zy4KNcabuL+r2bb8CUKoHyuTb9bjp0D8SyxW8I8V
kyxfqRx56pRpyrFJPitjvv3Jf9xvs/OiwSKGecPzTTTFDHht3vgrZZVgDoalgsC7NeiOdz0HucvK
kJBYhkPBnn9hO9OCGB+RaXdxfOsellamxFRJSQ642HNXqf2a4FsnXDjVA7Nc2jFquSuQfxqdxMDo
UU1/C/8XgSA1CnXZhznRbJTL1UVU21y98lM1rErIy5si3BAnW7TL43uhnxVv/MIjgtVxgaZ1Wlmz
IzigqSVee5kdooDLBv4p0qngBMzkIfQcIe2fPqlPlyQysQNdDuf6uAM3sL2GqL7izIjhfSJnzHm4
Jcf0Cgfx+1TwE9mrujcQc8UHkjC3/rNzY/i9kLw5RUS2kppvqt6WpBwLpzr+C/+mt8H1RmgSg7sq
8rVIar321bwA3tSjBSXFTa6GBDfzqCat3Dx/MgqF1s10SRlYWr1T2hRvCfRfXFPdtHma0pzWKIZ2
2+jUpJNAyHBwUWgqY2K4Thjysm/UYrHLevX9xOJdmBSc+nMa15I/1mBgZsOsQ2Fixi23oEXpF0ZT
qXHGY+2NGlTiM7/+JxEc6K5hyZiGRc2Qdl/nSEXer8QMYoGdAP/bCbAsINrea5dpuK91KVKnbTn0
AYzX5gkowHf+qIhSozExonqscH4jr4R44gO51DN5TSORr2Zzogq60Lm4ZwCgatnoGg52DSyp80Ri
f0dkBbZ0+/adW/Mad9/isRZ+Iyv4xZOSdMeZNQK6+OYCR7FqsuEdYOmugjnSFYW3JA8y6FrEk88J
mJtVMLrrJdB5xYLicZSeFtaQVwantjFYjvS1zmIHt+cWLdKxA8tGey0Xbf5q6AzeKOxOPAn5/ppV
QndiIGQF3fRAfERF3TuBUhPFKWn4p4Vr7uPY889IGu8tM3t2FtgXvBUTTPAhwrCeTxdpbirZERcz
ypjl8NSuRQoaH6JqzNmQ6eT2l2G81aRHcpQCKe8SYo0QW+7g8nDwr//3Tr/CDmpnoieCmv2LDDHc
tRPxnEIenO5KPsiufsfOt1cUJN7PIeGTjrDDrWLQgFx9u3gXZKdl2rapSY11EIPfyg5isjULcyVB
1EIxUCTVB2VDsut+QVWwDC5eNANCKJ5xVK09o7xEIJk0qbgnGkUh9hNu/BDptxP8bPq/u5cXb+qf
0noL81hmz3woB6hqb3BES86ZEh7Ms94naESo/zT2CWuTS3ykhWkOpyHUGPAFjh0660ZBIrD0/GD+
CBQQOsPhpcNPExQ+ph1YT4NcUMT/qhPPcEgiNedz11HvP6R3RLKerjF9t42wgqIiADN7itMdx217
NXQnrTS7SFrAEuyEhokd7biJwIwcGD0Fw3CYMbjcuDlPypxA1g+DmOQraCmkAqer7fjIKu4B9H0m
+9pXD43/xT0LR98bmLSiqTm2D9Qqra/lKTGg5VfFP632IngzdqTptdvnHps6U0IfJ5Ye3MUag6Wv
iCN4xDjwfmBlVHvApcqdasU03eTSVgASuXBEOJztK2116WOWxHnEM+O8cCd9e90gs4HewO0bv3vy
dnmYCzhzDnU1gGF1pozeQgJ6LYcDG7uMCmPU+D/nm0ezq0g4N8V09qw/58sTwFAUABIMI0c0kAcu
ixoagKnVGlPsvoDSYZzYXbfCiWyRBZbsMk6/OD6xZ1Rc+SJj9/DfmuLRWk0TixU5o3sh21BlWIh/
CzpeaWI256RFBzYCL40W+mE9uKMgePG8c3teTZhccbimbPk8xc6qLVjwX7SXwnBqUtLLuHiIU0u+
gF+7b1Ibf/uh/nbLF8RrO+v3sDwHFiD2Nn5rnDiJFLG8xHUvb6x91dRG88mb7Pd+/MfbzTCFZ2sm
W5SbuIyQcYWFrpsSRONrscQAn9yblo3wBVHoG7uqO7wtDYZJKlv6+2fwseS6fBsgax5fbNv4JBjz
K9xbg5eGFYbFPfXPrx8KazBETTDVS8OvZwMeLG9i65kojyEZZI3oyXtpE8uF5re6XJpKbZxAOZ4N
qxVG9gmDcDETDZ2jpUt9DSOVUWpxBCKvmi8gdFcMP3J+s1bSaIZXhEA+JxwBrikIwF+OkZWTr0B2
UVKohkOeLEbmN0b8d4XO0cNqC0rxg+yibQITIX2WkfVxMPUhXtOxa2rAz3UbzDl8jH3YIqHA5O9O
Hs+lY33nz+ooIAWLl62+VXrlWQ7CnbhaEh5PsXDSnxVVzt5TBz8XC0lfGzK92FZXmDsVzRBHmxVF
4pOrRK9/mverlwxb5W3Q11vS+3KTGUylitO6CMTgC4lKlD5Ufelee2Jm/YI4xtqg7OJf5xp54Z4I
hQYq114ABs+rel3ebrXkfkJtrrCboipEbsVNUVy0iQSzvCPOTxwUXSm3JWDTJwxUG+XCWCOBpVip
LUpZbYqVTJ7N6ibqFK20ZFEuvONZlkO/61T6ZhFlEMN9X2ClTiFmYCVfh7/XXw7vJrbAzSsU+AZt
DQ8mJEo5leAhcfCLTahfzrK8mj+jThChgqlk6VvLSXW0LO+QvatTBb+IYO97+eZ0G3J57WHtCbAE
rl3X+aykH7KjRYcYpR0Qp8bUCXH5UeK8n+x2mzYDcnXbuNnI9IUXqnQrMY7XTcQErrv8iuRb1AGZ
i3Ag7ezz1zG3vh+vwekVZyxmL44erOVxQtokOspKNig4b9b1kKux1dRzluS3y9h0KOzpqMtQZo6i
uOwXFiLy7ESpt2D6ciFKx8j7hfgs5affeY8bOHY3sxE+VeoyjpkSqub4ICVbs8vvUTa7i8yk6y1v
kJF9Xbf29Gh0N5sWl5TlYKzUs/JGgkFseb33Z+RXVz6mWZ10vrPXjPyT5P8XXUN3rtKjgmivGA9v
coorNQP0SLrQgyehcoibOYTA2cog5nrkl/3kl2fTzhdYrukdGkMnGyTFvJvJ689n/LAGnAgDfv/w
UuylqEVUq05RD9PIi/b0Seb56OnLb4ZpdcpPjYTExsKZCjrpu/2rhAe4odzKyvHl13GqstJDmcEi
xGKQd9dXWUdscuE1ijjkeRkWD5PpWiYq81N1Ud2PaptgizsvV6t+dHgabaIEEWe5BwNo7vRn0ied
IW0+zrL0NaMkfziDt+Fj25Yi/whnP05OYw66RPP9zzvsaGELOwseP64kzjN3+afgHXC0hjPpd/np
RWfJv9ttjVGSQZ8j88VfTnIXs8G8qsJY/gz9StjH0S83i4BIijir2zjE88z0BWYdrM9S+trAgo6t
SdFr3gARbdtTHLrcrH5McAHfu+IXbGJIVsLor3/4S2saljkEoVGDX345j0PGN/WXgK6GUxenJMLd
ooMMbZsHpfkpm3Z3K82tbChHTFSTHZYoQysAhJm/XaW3fOK62VEa871ftEBfxfbpQsnWHbYFUjeF
1ub2MZZnyrCtePgck7az60W4qtrP+DhM/3JeSLmq3cQONsc7rXf0l0xf6ZVaduWiugeCHj1NAiAv
8DXI1FRv79W8M1ZapNVQWLoNEWaEBZS9EMKpOIQfhzrhAh25Jwu2jaqz9dQa5UH34JV0wdFzGL7K
9QB61m0ou82MXMB5DWJ5VqYmw4in67CEr7EWTSw7VtgyxD9L/iCOFAWO2vi37oTsLiJ22FQo+8eU
ITuV/p7CuROI2Riltd6ufx2Cx8OdOz0hsZuyoJtMmeR3CtLe3Ml/B9rOwF40q/THvkY15quC2w4G
fDZc5vgGAsuxZyLHDZq1oXy0dklg5bFgSQZYVMHE3d4fWTnimpxfBiX06wxE/b10CNn+ru7h80QA
bSt9JdQeCtulZ/QbnYAEsVZz1uyThTJ0vOiAhzFZM89tIZjuBSpt26sNGc1DHbxmTWYTDQtKWUkz
VHPBFnyFmjqGqVNEYetHjH+Fi+S4A3sM7hV2CmQ/UUmwDNyaBePX7yQv7KYVE0CLg334fxWNCXJ7
ZC5guhJTY5+HZ1rkpQwQhJEpsZsvSf3hco4pdqgKSegSkyB7SVmRQTCEd3aFmPVVYvYdFoobAUwj
diMLnPeinReEPxT8lF3Mkjo7rRdbOcGJO5hU0fGtBSlfdXXTacF2STDHgwlXzJubfym2ThNbaMx0
+WUk7YsBYfP9k09eGuykiTBOjuQ/osPSlb9HGf8LC8qOGJ7Acg4ckV2OFKzZ4p/CWIIXnnS9OA5d
mWYIIu5m5Qu6riDddWQ3YwNf1zhaeJ+7mraZSBC4ZNubFm9Aoe6sfJNpw7NCAcHPr5E2voOjLd1c
tvRtRV7zDK3VCiwhSJOk+cy9XMzy2dB/s6DlGaF4atzID3AsOl4sGRbz3VYiWPyottW5XalHx/nu
uFkpGWvVbtWJuW3hfIj8mgcxCV0cE5xni4UdVtb76c062UhI7lAIJTe6QMlOLU2LP2MXUAjIDSzh
vV2Pc05nWY5sIGvwacrumtgA1S2rWNfVto5UDY2mkqocYjYCoUvfNeFZ7JY0lFytS4sZfX3wNVIC
0TWpp4+JH8Z8uQ5gWQe8Qj+ijGJ9l8oCUs6Vpi10CwU5hy0fqI4aaJU+Hpqu5/V3O8ETn0j8cOMG
YxjboAAVo31J2AYkGLBk3ZZp2hSH1ZPFhDP1ElOmdUI35hVE5NQGvQATrRheu9p98ViFJbywmDuF
alwT4/cDP4BAV7gG05BYq6H7iRtiTEMJYriLJEzbAOR65nJ93e1Ar1DUfsuvbBuTIKXkSLuCcJP3
5XIpgOnlNuq50HKYNKZ5RWK9MODsVZbdo2q+CYhAp735sBqxdYvn+B6tpbAHqrBECEdoCcJ7VSJH
Zw38GNtk0wTk3HWWQf0QO+C420Kalg/9lYjwO/12tiSu8b8Y8FPYzHBUqHNNX3p0ugwb0MEt7eFF
2LCBs7O1TXplblFTrdiFBII3LUkbs7i8p/oxGhpU62KXRPZ4xmR91mATQvhrbiNg3HXEWWejckRh
ztslQfE88sQRyXZOi5+R0bSZdj/clDlM42JmUFE3Q1Kcd6fIzFGRpV7P5xcg4vDkICi3JkFgt8G0
7F4FAu4S2QwJP1AAAxL8zDGQjjHrp5SbmxoSA+b6txSkkIVpOGf5/VfAFefMTqRBhEyoCRc+a3tB
i3jGNbZqVXvn+iNN+Q0V0Jg0A48p4E1lhLX2DnmoJ0XPWUrK1vDqO2DYV1wZLRNHgaPMPh8etTkn
3nPAkBDYV1yt6DGo598fn0jHz/FzpjhU+hCedWXlHr3/BhjiFXm+BekBNad3qduWz3B2VwpK0Q==
`protect end_protected
