��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��,�y�}�ǰ�=4d�H���`I"��W�`r���T:tB�T4D�m�)�	1��I�t��
��8(�8t>s)ו�."[�漆���]�~�]��;�O(1#5���D���d3�q	��9/�I�w`W?ދ�S"K7��5�,l��C���
@E=D��!
����荾Z�V�h��c,Dt��&�����]4w9K_9O�=l�uE�w����[R�\�zÚ�-J�$����åCj�[�
����T=���K���h�����,������#�z~��?�G���B�~֨1)��k��yq�$/ju�YA9��SX�{@��mWt������w�F��r���������O)�mC�&�����$��^_��|�����=������A���_"�s���50��-�ݡ��kVE~�cu��'Ah%�����v2ݲK:|�g���7/��=Q�u�~��qC���
qSa�a�n�m(�]�h-�FK�]�Z<��K�b�s��'�����C$Yכֿ��h|�[@lXJ�*Qm?�аR��(�v�vlr�j)ڦ��0p�s�bv��jy�-����(��N�vהS��Y�n)!��\|9��;#�o:�#��9|TWL��L2=�'���$ƫ���19�?�:H�A���T秧���,rJ$�p}�a�ڡ�rn#9���~�1e�[e���!������{�T�7���O�z�������쉎�<o�j��D�7��lS�ƃ���F�V�:¦?�,�:4I~P�o6����2
�ԫ�#��G롔�qH���'> x������>I�nN1.�yφ�V�ǹW�)��	�3���k��c�Rw�buRA�8����\��L+p����rw3v�FF��8��Y��8p��s3jL&���9>��y�(9=���a��;(�AR�cAw
S��k+o���⋠'O	�iYҤa;L��g�=����*҃��aW��@o���:pÂn�'˦N!8���%�I��E/�;�3т�v�n�.�e�B�z"�Ӆ���z��6�G?b�9��Z�Лkb\�)�s[X�dp�_����< Z�׊,���:k9��� l
�?)Ʃ��,�E�4���2����c���#����\b�u����x��q���M�V\�����/�@��Æ���C�)��N1 ԉ����V"�L�z�%e�й2UG������{���4l<h�`���}����pUo��&�eeq^�i�1�lz�Ղ�>��*=� l�Ǩ����l ��<bI5ȃ:�c�y��@
�K�y�~�� ���H(M�0�w�-$=��u榑?���8m=`S��I��v_�#&-QԎwo����&һF�A���|<��<�����\��~���p����Q����ݹ-B��X1Ɓa��ˑ��d�{|��
�	g���v碄�d��X�?1�pEKֽ�d�݇ˏ�M�j|��0F�����N�&,+����	�q9����| �{���Ҫ��hX��_������푿����5o"������/F�s;{ɛx�^�WU6�L:���=��pE�2�,~H�|����s6���_3��?�1�H��G��ʼŷ1 ��M�j-�g�QP�,�  n�P���??�������FO�pn>kgz-����f���Rx�0��`
2����N�K6n�;� 6Mt���ګ)=G�ii7�Oq-)�.\��ߟ*)��dL�ȍ4t��rܳy_N4�˘���X�zGC%޿�]gcu�?��y���.'�?���l����^��^���fyH;� 7�qL~�����)S-�E#:��nh��+�8ť*W���N&����)e|>��Ts{Ʊ�5���/���1@3��k�d����D'��!�%������`������-Yf�8��"O��w) `�5���A)d;�s�k=���Ï^�t���G���I��8��1�e����ݿ�
EX��o9wuq� �^0Z�D�Y�$sB�0�Wj$!/$�h��g��Lȗl&h�'���[�����g��,	�͡��اe�YI�����4�_��z@��5�~� �q�D��[��d����!���hx����q��r�G�k	Ѱ��5~��hߋ_ߌ�����C��H
�A���F)��%~��� (�%.����X�˒qL�[�jAֹI�eT߭_�.Ik��9p5#���4��jS|���d��o�ŉ, #��&?`,Aή�kM�LM��������"��u�z1���1q��I�%��^����2���$$���^���}�� n��.��HeTuE8S�ȓ�E^�-PA����4�a�dV���t�Xʂ��fp�uD�i�@�v0}u��s��ٕ���w	��z���Y�g��D�QMs�0
]��©̶_���d"r�L�1����G�I`|J{�7	
G�!�9#�(��\.b�t�^����;�O4@���6&}?R�>��w��c��a�G���@�ӟ�}A@���U��u��w~y�������C{98F�#��w\�{e�ɫM�f�����aV[D>��	nG�j3w�9P%HK��AU�T�%!ø��T6���6��q���X˳�f	��^�c��l���E�n����n���7��l�r���W�`oL���""��Z_�9WƔQ{'�)���	d�Yx�.<v�ڒ1�v�����������;
���@{[$R����#yYޯt�%�uM�g��.�ݻj�p:���0�����D?�:'��.�	�3�>���@��\����F_I�Dvթ��6h7=q�pt5"�/��Υ�YaE���m�H?�Oht�S�q���]75�3r7N�h]��s�P�:Q0-I��m��V�>4�F)�d�c�F�Ӭt<9���l<�á����~+��G�x��Ȭ>_��nmAkcf�ůƢ0�p�*��=���.o�͚Uggs�6��u��΄�m�,��I�uq��^8LOO�1�T�����j>�
�F^H\<�������6�>�Д	>�p�!�c�-XB<��<%��`���d��mO��z��'�@����U�G���GV���$�� ��x���Jz�;��F��Ş=��R���3e�!��E��X�ku�N g�p
풛��H*u�>������D[iܮn0w�<rp�� a�����@�^�������fH�Z�M}Qbp���Q����R����{�b�m[��iAp���@>��P�#Q@�*b
�x$���f^&�C��p<9�zl4�-�GWr�;I�#Ez��n�I�۷L='�"$�1	e[�M=)����8��<5������`�^��[6G&9~�H��<����\����{�z�6b7�#��ɚ�0]�5&�g^�Ӆ�Q�n�@��gAe�Q��G#���Y6Y�{�'�4DFw�T��Q��OQ�ܓ=k�9��U�y���e���.��X��R{mЗ������f0�|w��.����(�`��mQ���4���s��`��~�JX�>19�S��v6���э�����5�����2\���<�_2'N�|3���x%Ǽ�'�W}z7���W���'��� �NE���R�y$YH/�p��R.�9�����ݬp��0��,�)�5ɩ_J2#d�1�����@IѼ]>)׺H�ǒ�'k7	�s�8�$����7�x��6?�u�<߅׳;0�>yN�׳BĻͷ�9��g�@�l��tI�X�K*־�{� �jY8l�����]/�|Y��^�/��GM[���yu��@T�!#�v,j�fL�H.��HED�\ƒ��u�}|�L�
Ak�
�&���y)���ڞ�bn���b���f]'�n\~G�)<?�wϡ�P�f�|1�2��4B�an�+�)U�҅�Q3^���318�ݻ'��x�����?����ye�"��JKk��>�v�RS�7�0��}a�b����b
��{[U��^	a��)Fd�:R�|Pb�0`"N��2��>ԆH>~D��k�d����y�������/�)g|�,k���sv�4�����I�rN�i~(�|E�K�B�����A
ըD5���?�g��a-{��U��sĦ=�I.ȤV.�Orݬ�!�������0p��Ђ"�{�?������4���"����?�W��o�HE��!�x◮�CHY���bx8���c#5P���H�"U�����kJ5;�+��mz�����<�؉���S�:�;�Y�E��\��m�p`�@Qv�2I���|F��Е���cE�7��׸��ס6f:;�pξ^��8�PP& x5���2�s�'�s������ap"���ݠ5�UT�T�Z�!/�.sX�U8�*҈��*&��H�|��er2�c}�yL�]؊N���<��N;A�B�f�l<]Bh[�m˸�mʛ 	�khC�N�m�c݂��Q�E�.����Y�<�H~�f���g)<%~�qI��jzŀ������ىه `̦��
�|�����l�#���jY�"����$����C�m@�5)�pN�-������cy� 6?@�DW��q@�ٽ�s�&41�ӣ,���G<Sģ��6�N���~�g��DI�J��]�-�ͽE�RK���G&��E߮�	(���f��w�1�Y�{r��I�z\�le��_�5�v��0�ӏ��|�c�7W�@���(�T����Mɡ�g0�?fcQo�K�������1G;M��T�7Y���)�����/����?�5T��ݘ�f�Sp/�kܐ��zE�1��:�Ja̬�W�+�x�M~ͭ��ZȌ{���L��1���5`@^�<W�~�֫#���H`���si>5\�Zǉ#}y�:m�����N$4?���"U�ɕ��3g�_k�-��uU9��Đ�W\[W�i��E5z�Ծ�5��h�Q�8+I��b���D�8�μK\��bc�X�pM~�O�>�,��Y_"?���*�2dB{"v�!������`wH�y���F����w�;�~Uk>d&����������"=�qX����@�P5�T��_JA�n�.!��931j��F�0Q���=pOk��0�Ϲ���_F��D�M �+�2їٵ�	eq�Z>-?��j'0j�h�EP�=�wĐ��l*4�T$J%�v���1�6��FI�;.��H�A��&���=s��hI2�E"��uck�a%�3�NL6n]ٜ����c�����PruO��bt��X2~d�و7����|@��r��{�{�����F��ڀ�^��>
%K��EUk�)ȥdڟ��y�yǡ���嚻j��s�dx���m�H���A'*Q�_dp��w���ޱR�	��~���6C���&%<��	t.k��a��1��/x���e��,��.MKM��k���'M�9��̲�����B\�rQ��l[Q*�����~j�͂߃�'�k�XbK�8V�ڲ�8��s���LE$)+��˧��_��xR��3$-��T�W�@9���[�r9���C��Hě�ٓJ�Ngd��:]�i���m/8��z\���
���o��WE���� F��ݣ�dh����-A�����7�Mr��Fn�Ƶ��;?��4���^{V':	&v��\�p�K_�<h)׻�%�-�j��霼�{���-ߩ�C�#�(b�1n�eV׽N�Xg��'����F�|ֳ
�(S�����K�1�S^� D���%ޒ�Rc��C% �Rq�C�q�
-���K�*
E�Q~�c�5�&��r�k��IB�nzu�-p8pK�{�hV��8�~��T�B �Μ�� �b=MUBH#�}�E"�d�tV�mgO-��~��`���0�32�n$��F��;Y��Ӈ�|�#۽{��[e`��h�Q�h[��0�W2�H�R�.�{�"���,56Y����*p%~�=�	��͐9���ΏA���@�Er "h&nP�J 9/ߩ��tM-eMyQ�&&6j�(0�����ӓ:�|�{t����s=�k�$��B���q��i9�5Z������co�^�f�<E��#�deU�VŢz:NZ�}�.�`J��6���IГ��.�d��?Ϥ�aY�..�1)(�[n��[�йkE
�g���В�)ee�>k���Mo1�ԫ�����q-`0�[�0:��:�:̎��k�6�O��;���S��(!�`EE#��3��hYW�P��W�Z��`*�g���
�:R|��a�D�7��8�0���P���ʶ#��oa��Zf��6H�fҫUʆ�/Uv}����A�}��BȾOo5� p�g��Dm.�<�y��������T�u@w�/P��x+�i4ȭ��0�찵n5�I�ꀳY�U�]�-l=�(��g��搧��H{�W���	�3-�\S	�>f��}���,s?�{t�#���K��W9G(���zv̙r��J��N�8��v�rM�ٷI�7���pa0�>���f��1��uO��L�$�ANՅOɉ�5�V�+ݝ�!3^�Tp0.:�J}���$
��zw�L���{��\tGEH�� e:�֐���C�����1[!�xi2���gtŤƻ�2�!��]ӳ��P�HH~�T�����/�ԟ+��`���;*%��_r��h�j������!������!e*̩����V.�9�8����RB֍hdʼ�_L����R�� b��$0�%��7q�T�r$|��H^��1�KB��Eo��ЁT����9>��Փ{�ϙ{�ɌCfY潡Щ\)�݉]:v�ߕP�bߩޫ+JןR0,�o���+�����'�h��M���K	�_l?�없+���<56=���cs� D)��O���k�TUQ�!a"��dl�jdP�y5�������}�2�o�����-��q�ON=-[����1�:pTFK$���cP�(a��yɅ ]TĂ	b����	0Ȯ,ywq�𵍗?����"���)���$a7�P��&���D/��*������t����ek�Am׏y�L�%g�e�Lч�'x���?����~����0�m�j�h�%F�,�zb�R��i!�LT�S=# �[��ߪ���2l(��� J�h���c�X���\�/��d��!�&_�D#��	n��^�o��S/~�]�w����珆�*�g'�3���*9�9a��R7H(="f��DL�?d��Ht��{A6���o��B��8�c��z�&�hW���>~�d�-���BИ~���D$�!z׭�d�%�V�U�CZQZ)���)fY	�:���	MSaxX<�����{s6�Mf\�O����C
Hݬ_�0s\.���|d��͆$t躟k���j@5�HS�!�qi�K��)c�DQ�#��8�鰃��:�n Ln���1�UE;��o��=²�Tir�@o鳒���#�L���2�y������7�R�Z��Z�BP*2�S��[jv*�ُ� �c)�R7;�3��p�"q��lb��p�Lc<��Ūm��R�!��q����ő�
�Ts�U8.V4{�e��ZU��}L��'���=9��g�K-8� �l����EŚY
�Mo�`&��/�?�����Cc��N���E�0
\ֻ;�"�њ6O�@����#Psȃ&k�x�g� ��]6�>J�G��m��N�l]>��.od2>�̧�*�{Ǐ�$�ѰmXD�/i�,���G)��|ҁ�y�ǂ�yE��1�~��ŧ��SHA�ߘO�Q�.��Q��*���p�^�-�c/.�;��Ƥ��
8�@7��l��][lg�BuϏ�����m����^�aK-5�i|���'���5RC�3T���79	^d/��T�qT�Z���aX��t?�~x2�,җ?G^�̀��c��w7��7x]&�.?��ً8��Ҵ��
X��r�;������_T���
w�o(
F�w��V&x1��JI� ���N�F���#�)�ż��	���{�<�MJ��mmy����fQjT���+����{��ȭ�O�!|5�h.{��/�?��L�@B��U�`%���F�����3�.�����;�r�*��Y	�^ѓ�Fr}>g����}��v�y��ہ��Z�֊���7p����V�� �!�1�܇����2��p��یG��d����@�,��0V���n�ݓ���6x̮5I�������%HF
W4&�qP���Ʀ�?�r!_7�`����O@�X� ��jr1],1�*SyN�&Q�u��-�ݨ�٬W���~�V�Iv��-�>z�ySX��\���F�&�����܌�j�#bMJ���dA��
��D����9���Dv9���H�����m���Ѳc�]�I�TFJ�{�T�����M�?1�=i�K���q�6�2��<�8ZC�>Ȫ]�ij>���r���t�*$g�s�p�ll�8�ХT��&�+�{��h�DB�l��SI�����$��K�DK�<�XK������n��K����9a����(�Az�h+�ķBg�O�<~����G��*
�)v��<�u-�#�]%��R�H�Uԙ1{���P�/j�+�\�v1�s��0�ѡ����f��sK�V� ֘s�5o�����X�\��FX��^6���s3+6]�"s�D����p�w�ϫ~̓�����&�.�j�M�W���4�#�^t��m+���Ox ��^QY����������սY>�Ӑ+�"�k�}�|��T�:)���L��~��"�p�*t!_A�K�]�m���T�Ү�M�s3��''���|tΔ�V��fq�m��ϑ�mV("mS�x K>���<?ҿ�a�����b�w��"4!���o�	�w��R�"��g�F��,h7 q�XmTv9���85���<5���)^�
n�̓��[w��-�#�d���Nׯ膠W.�U������>�����8�"t6����C����b�*j4y�%Ur��y��=�fx��Z�8��$}�RV��IRڼ���.m��.�n�f,q�& M�jO�<L�Ԅ�U�F��^����3�N�CY���6�Z�����ʌɿ*;���9����З��(^ړ���`�8U�C? ��.�2̑�aU�s����#&��R錅MyG �|mjzS��=o]�!�m|���"�ֆ�?��ۤ��,ꓫ��<3'h���瑺-����=�|i�ܭS
����Z���R
i�CR0���,�uI(P آ��c�~#�g��X���3���X� 6�-o�I��k{�I�a��҈y��֤N�S�A��N(i�.�zSv�`nc���Ul������͂�xK��$L�A}�4�7��S��l��@���o��*�m�s)�|�N��\��.��?��'�w�H�w��b�=q�V�5�AyY%�b���g���3�<M�5!��(p��{.���7l�3��u�%4����dT�͡o���S�>��M����7\!�V�����<EK���c���}���޾z�����~����u��s��FO�)e|!ѣz��BlBb8T�_0>���=��4��k ~��Ъ�(��@9}R��6o���|��*��;����I��o�=�`�B��{�����|�<��Q̘E섆j��p�/|&5~D�K���8���4�I8㘱*�n������P�h��������X�gd�?�O�~ml����<����QsFfQ�v*���~�Û�ǭ�N��(���J�f��I<M�5�6@�'��6Y-p���O���L��o3�;�m%o5Nҥ��)��t���J��kvX7�_�K8��D�Fw�Ķ�p=��f*�|Y�{���'�AGI�-w��_c����R�B�vP�"�c8YV'ɧG�c/���A��;39hN� �_~�B�"9�e�	e.W%s��1�C���<�Gv���\>D�7�Ri�	���8L��:�lq,�FV����D��Qfe�}?�S |-9s�&m��sV��ܞ��|���(M�[	���|Jf��=��}���[�p:��z��ZC}Z7*����S���*��S{SoWU_�Aq\-����E߷*i��+X�(�����52�c$x�7���/�S�rK�-J�"U.�>I"~s�W�.]���h*��/�@'&�M�d ��c���(ss
��V:;<�.0�04����p\Sc�w�v����x�g/�wh�_Ɵ:�ZCH�3���T�_�]�bZ�l�M�2��v��"y��SET����maf6�E���m�/M��E�\iX2+R��(Xg���w7ph�9��u�D�ژ�Zf�;����zSIDZ|��B"�`��J���]��8G;�������C����Eӱ�q=�����}Ēot1��,�zsH �t�6q;�le��� �j�E@Ol�TZ��M*�.s���w�l��Q��͟B{
j<�����MҸ`H�d[77�xt3�rĎ�"��cS��a�����0��c���JC*��7H�Hu�9:�5b�0��,!��u��y����B��S�̓Ϫ{ks���ݖH�N�W7�9F�����NΗ�}	
R����wY�AAM��������O�q�i�q�Y�R\���O^3���]6�,����]찈�k/��Aj[٭|��n�z�����M�j����vW�Q��F@���^����I��G��Q�4_�B�fȳGQ�7��&�=|ǯҮ.��3B'�,��a�B��)�q��!s���Y3�:r��(�w���4�A-�W9�b���*s��F0	|+H�U6�Eiz�0���;ͲUș�~���Ql+!�����Prmh�'�����?�r+�������,*I,ZK��a$/i�̠R!R�����1d떵������;��6e�Zy��Ѱ�}T@��3d�l��D���b��{���.K�����(��?�G���N�S���fi�)2<����h��snf�[��b���"�=���v��jbC�{�X#p�k�CK~�G�WҤpd'��9�x�r����S���pAf����:[����)bc0�.���6�z���}���7��׳R�֤�<������ք���;4f�~��9�@1�*}���Y`D�,7�{d��s�۾�A0?�T�� �<:sO��q}+���K�t]�����67hnyQI�&�}�AG����r�(p�ʑ�׉�C�:�5��##���XH�P��"�s"�)8Q���gKKi���Y���[6�&qY�J2zQ:&�*��'�^O��[�o�tq$��V�;[��.�9�h[�`��>����Ec�!sM�qC�t̴,t��HMM�;�4
a�W�E۔����02��lR�Ue�h��#vc6��1ͮ�6a߲sNR������#e�0^\��F��Z�ܒػQl����e�B����=��/�0��i��9��@��8���7�\���$F��e���*`:�� �e���zM�6uzU&����<a2��O�/vZ���y3���� =g:����L��!a�ڴ�q���k[ȡG��#�#��L��M�,܀�~�v+��{��DT�}���A�eT��k�f��8È�۟�'	c���+'�d�������wH@����Ύ5�^�t�^��`�/���B��mTh'7�X`����.�v�	��a�u����v�%x"Q�E#W���ro~@n���=�kw��t�5�?���"*�Cu�I�.ST����c�6Ϳ������p	ύ7�����E��yx;����u0�%P���<���i�5B��
阛X�V]�M(�6l��į�Q4ƥN�I��$�-*�/��&���-u�t��- ZD<���H�4\61�ؿőR�ļK<SpH'[r	�]'�҈]�	ta���|����r���ͻ�ęA,����p�D1>C�bj���!��ͣy2��:~/M{ r��F�hsӅ���*�aX��je�2O��Yk �=��ֱN��\�ˢ���in�4�&�0��Q.z񋖶>v=pZ��8B�W�?�}���P���k��.��
����~�*QP���_!���+�)�~�؁	��'3�*��z���J���a�x�S���J��i��J�H����$ʘɳ!���E�Ż'��PoD��w��/Y�d'��z����Z�t?n3��s��ɵ�;�_�MW;V
�Z-\R�5��x��{�~�I�+[�4���6AF��=?��&^Ӆ�D=�<�4�c���ex� ����,��/�啚�0f�[�J��n�nn"�n/K\.&l/�^�.�D�[7���-i�ެ�8���hR��E;�(������4b�}�&��&�}��ignɲ�IÞ�����N��nk��ؙ�b�@w����?�d�p6Fty0�H���E�|�!�ݞo�}�������F��(�����R��H!�7V}�����,��4��c���b������ }��9�&�Rg���pC>O�K�r�./�zB
c��C�VFЬ��ny�T*�	6}���5��<g���wp�E��0f�V�T�>2)B�b�z�Cߧ��+����w^n����l����O��}g�.����5剽����u��R�xw�9uk!��3�J*O�����Y1�5�T��V��f����'_\Q�D�Ht����"Ι��l	�r��y`ϱ7E3��*�b���4O�3��,�𢈟��~�|�E(���V)�X)}������3a`b��q,������.��̉)�v�'fhxHċHԣ@��f������$�,~<�|Ү�0�����<��z�p��2��)�𑵢�0�s!���8�+9g�'�8ٌ�����^�sR[ґ����2I�n3B��5d9��{�uG�������� 3kBAe?�N}_�Y�Fz�0(�JQa��Z@�)A/3P�������؊^|��W��!���+7�jP9�` �+�0�[�"������J޷nJ�f�TMS�	��TY��G�*ϗܵ����gƚ��=2Y���m׾'���Ƙ�c����;���s�u�
�:��Z��l��8��Be�8ɾ�$ۗ��?�11O�ۻ�QNvh���M�MI7�ZK�;Vs�h�ˁ���u;.x���S6��i����ļ`|����5j��z�K�k~�ZN���Zc�kp	��pM��BRl��ӈ���E�jw������KRq��,��ɝw)hZ�V
�Hmu"@EHM����b���/KL��,É7A�Y6
0����Ax���s*�Q=�h.9�+F*knT�G�Qc�y/��
ڡo�b�e���1rj��rW�g��ߨIҹ���ri[]78�K����O5���+�띡Ӳ�_�GD#PZjq,�R���,dfV�,񬩀�y����?�jQ�@.]��w�:{�$�ݚ-u[-7L0���`|��qG�*[Z��x/@2�c/? �l],�Kfc�%Ɔ��$��ٗ�9��k����2
�>X���%go }\_D��2�U6��pH�)�1;��Ş�����-"z�Bm�0��D�5,ݵx������X�Y��2��e���;\�#�r��~Q�\�ӟg��-�+k%N�=�2���*$���]}1�ʕ&�ub�׈z������$����Y�m9}c<��P�\�8�W�vO�9Q�fV�٧A[[S&r���e'���.�h�b�ş�-N���j5��4����Q�(�џb|���T�� �UW�m@W�B�i��e�1�2n�6؜u���[��~k�0�����1�P-��q����~��g��ī�N[�w��Vq��q�x��CN�g����pJ ��{����:k�7��o�	3r�=�X�j��A��e>���ao�>��ʷ"�{����:��P��r�2�>�&�F�WO�W�]Qi��5��O#�W���-QE׃���&GX�C�_t�
@e��d�\%є%�il��Qh�K�T@a���٪<\�#�ß�lZ�hTx��YA��H����Ð��
FR��u8W�Z��#)���Jx��-����L�l�����%?�Id��	�O6�f��Ov�@	�i2jD2��Y��8`��fF~ڼ����d���ߞ/�+
��� l��avYЛ(����or]����	�s��\��G5�c{:R�yŊ�C&�'g�|l���E���;�m�$���v"n�XZ�ZG�����7ȑ�g����}Ƕ�����Ǔ�ֈ����4$�����fGH�����}���M	�mA3p��$�\�ړ��p�
:�.@=�*L5���I��@%�|d'�5�9&ڸ��'Z�p�Q��"��H���c�X�g���A��t���*�3 ŴI�m�����]?/��G/�������\8��ˊ�b����v˴��A��+oQ�~%[�\K�D5�4!�3�ͽ,uM�AV��|�)��t
VR3K�!v��*Q��b`���_\R�o�X$U�̍����UU���{M������}W��)�<]�gC��l�|	MVz!?bc�7����}l�G�#��G�IUˆܘ��u�Q�`Ϣk='�Ec��i7�����b̋���69�?+�(��T�({�@����k<S��B��o�TV�H�˧h��,\)�fm}�}�q_��0��a:�5؊����WE���z$�@�Jp�^+6����g��އt�}�ˍ� S��S��U���nC'��Be��`x������4�&a�/��x<��+^-e�A�aI.�b��Tf2�@�YFVh�_SU��R��s9>�2�=
+�������X_cA�6��F�Q��U��Gv�(@[l�ޱ.�<upQ5���0M_	�Mɞ���8�m��;��.-̈�ʙ��b������Ft���-�-�/��߼G;�wl̴^X.+��Y[�l���d$���%Ż:&�I!�f"��S�-�?��WCE���BL
��N9����T�#U�?=��HȰK�T��Q�q-��7����z���q�!�{�<Мd�I�K�����t�O鯸��i9hL���I�Y�h8��.��}]Ӂ8�B�٬(����	��T����B��w)pD��M�G����@7�[sY�Eļ�Cn�W����x���x�KČ�V����,x�f�
���î˛���z$u�	/�ݣ��;v,��Uz2�$z6:��r~A�w6B~�^��� ���픴d�4}N�~?��<[QƵ
�	�ji�$@	�r� z�m��#B�?1�U��2�#l�qXj�\����?/��v�.��H�����[�Ç/���i���M���	�984�
�e��8�� �(�.��s�d����c�'�ӃF>���.
�wjw�z��p�&oi��������b�pd��+{����G���G{j���r�We5�[��9"�*KE�>�C��NJA�	t@���E��CRyR^��;�+��}�2����	r�jŵ��r������fY�r�)=e���8E^�Oc�0u���dX,��Ϡe�9pδ͘q�U�]���Bj��%�D�x��*�ǋ��M���#�����^��ũ����LBV�y�{�;�%��ه	�) l���wM�h�3��ׇAL��pE���l�"��k Q��b�ίFB2:r[`4{�S琊tSO	Q�t�ÝTݯ;yߍ�qs���2h��J�(L_�&�?p)�+�@��	�/�2"|f�ۗ0�w��Õ-^�bY���l�	����)~��]`o��Nʜ.�~_���Oɴ�O.6�0�`��~ ���w��g}�Rxl�T���a�ލ�<����2���F�t��C��}v� �8���HmභdN���}�j������ִp��#g�=ڰҷ*���h�6g㘙y�����W��/�Cu�Q��%d�<ם�Ꮤ��=���۲Jx>�:ڽ�E�-�' ,ĔM�P/��>(�k�h��k(m�WԚa+;�
k.�*wR例�P����-P���:,`�\��=�`	<�0�1m�tn�~��.���~�6�"��p�ӳ�,�j&�_qG��z��_�T��c?����������:�aL�w���Tj�`rY �!RZ�����G��;�sү�$Hi8�d\��H�LSehv��R���;���7�9�S�ݓ��_i��,7�/&���4��G	�oip� ?������h�u��w���.��=�(���T��N/��:R���=�1���uY��ܾ�XK-�^>
��԰F�{7�?���Ӧ;��M���΂�;dK�||���ſd��E�k  Z�I��8���4���(�4�wr=�s��D<� J@[$��] ܭ3\���&�?�������G�x�4�q�V��|f��_��d#@kd�/Bz?�+���5��{���b��~��;�ϖ��o��ڡ���_��p{K���R@����UwM����ꨐVd&�`��'/Lb�?j7����O�L�Ѩt�A�B��9�<�4]� C��+�U!JC�N�~�s[ w6dӺ#�-Φ+�2ɝ�G�'mx��9U���E�C��U������=�qx �G��&q2?2��؉�,���L{�_��Hˋ�t޷x���8�?y���F��*�rr�5�0t]�[)��͒���`O�*� �ܼ�yw�=�U�(}�v�a���V\� &���z�M}#���-
�NgJ2�)c����m�+�A�a'�>��x<���~��k���cT��w��!��i�?xFa�8&� ��0&������rV�w=Kv�'���ʲL�"*{Ve?C���c��]%��j,ĩ5p	e��c��7��j��"8L P�W�W%x�9����NRx�C��#�����Q���1���I@�6k��H(+b'Q��O-Z*��2Y�0-9X2�xH���'V��Cj���	D�X*e�H���pry&dP�#�e'�]/ا�LA 2u�_�>C>�0�Y5c�4�d����#Z��i�z77�n9��R_W]j#wE2|'����Ydc��w2tl9�D��.�e?>8�!���Lbc�um����V��G�v�*cSD���f���pE�Xؗ�YR�eO�rK������L��41�`ɸ�F�j��2���q�� T��u�Z��/�V˔* d�����@��V&`�v���'�M��kN}њg�!G੩��e������|��8��D�o��N�-��?��l�"�2����)El+��8���8��s%�{b�w�ﵙ�7��L���~�yC:'h��+uJ��%�x)��|TVc���}�C�#j<r���q��Z*D��=�-��O�_���������`��bv"�h��K��#��*��  ��⿺�Qt�\<A��,U���}�V$)�h�nj/'2�x�SR�#X�����Y����P�D�U� ������%�=�}:ʴ,��2���f��I���`#��� ���c��Yqס�3��I����r��̀���O�����8�,i|���qi,�Ԟ��G;�j�bk�66`Gf�޶y4���n����o����toeֿ.-;�zhU@�I�=}�!k)�v�Za���.�72lڙ�n�R�㹡��'zc�"#�I��:6�G- �O0����Cs`9I��4C��Ӹgz�\���������S�D�
=�d#���z�q�
a]q�S�"���2}姛/�0c��kԿ-��#)覑ݰhݣؗ��6O:рsN�c���8'����|�������n�	�}餑ʃ����Z�	�����V��o}�{p��nJ�'�����Lq���0�[���k����*
[�O��D��wǄʨ�,Wzuj]/��,|=і\�[�XTu�n6��X���٪����y͙J�-���/hz����i�]�e�^��X}��F��#0�������%��Im�NDv�D����AE�
)��U�4����z��'�*��6�򆜀]�+M ('�/&ອ�;��S`���=~�A�'�!��ܝ*�
��Lpj�_����g�@SC�N�a=�cv�Fak���
߾�	#O5{����E��X�\VZe���;���n+W���X7�ף��"ǵ{���F��Y�R�!E?k�4ڧ4�C�F#ܔ5+ani��߂�9񷦃4O2L��!�����*
��פֿ��h��Ja�ܵ�ÄXH�5���v�H`���W���cD. �P)�ޗ78��zT�%�w��2�G8��o��{���urW��ƃ=�67�i�н�����+��"�L�돂ˑ����`��~�&5�5t�`�¬$�VY�4/�@��AE
�+(�|k�fx�b~sV�w�w$~�8�ٽ�\<jz���0o��iOmA�F��P-��e��ג�[-˚�4793b�}�v&N5�F�%	�����>��ƊX+�]/Z��vF9pC&�#��j�c{��p���4�ן̓d��gY�f�^Y>�����	�|�vf�x��8�RT���M�3l>pf6���A\��Cӫ���i��Ʊ^�r�U<��W#J���@G_��ʟ�0xR�����*��g�w�_��c�ƈ�$����6;�g�~�0E����`��'��K�h|A�0AD}`HY��/�+Rzmy���Sj��#5�2�)5��æ��1����@F)ejo��Y�MK�v��V]2�:n��J��N�N=����N��m��W�"��z��Я��1V��~�Z{Rs���
/���U��#��OJ�.�ۗ ɿ�Q�}J����dL��2(��9���-9}��	0��뚒�E������[Pء�dhSj�?�"o�k_�:���N�uӋ�F�VӇM^7��M
���W�^}9ĹR����Ԍ�� 	�b�K� ��+Ο�0l}d�U���`>�(�5�v\'�`�'rTJK�<�����g G�z[g��My�#� hL��pRZZ��jt0��
��-Zklp���W��t*5j�Xn�ݫ�f��^rw�ugɮ�T.ǅ%q�(y���}jت��Ҝ.���|h�����3��(��*�mf�x8�g("p�4�{S`V8djͲ�ְ&��D��<�4�3<�*��[L߮gUY1W%��A�����)l�G�B��5~�*�=$<C��;l7$>Sj�j7��{3�����o�H?Xw��PA!Dq��A�8���I�"��_ʛ�!����g��fS��i.}�ֱ�&�]��\��_���3�m��K]-�Νϗ��;&ꒊ��{�!jjZs�+&=tl ����@*~��f�d�pz���[�D�y�9߯9����N��E���{-ُ�;d����h�{���/��D�M��n�1p$��x�j=s�\^G�!�b�}�"S������	���q��E�?t����.g���h��Z�p��)%�J�x�"��?&@fE����X�0��l�}�!9�R����A�R���f�Er|ӄ ̓��G����a(n�{w�v��,2ٸ-^����̚dǅ��U"�Fٶ����<���-w�3�d�Q���%�x��ի��%����>��X���7XX����Du�w����E���&oׁb���ˮM:W�I�vV�<$�&���4�j8C��l *�V�|�	%`'�tɹ�|)�� Y��a�I>�H-f`A
���V�d����n�+1��w�X���U�b8���3 ��K,W�:z��S� �����vaF���3��KG�*��%G���ö��(L������5 W�Q����;��3Y�@L��/O���,<�~`���~x����@�(�[_R>)�� �&3`�xﻯc�-U��Cʌ������&`�(�?d�tT-�1�X�
�KR>?�m-z�'�h�#�b� =Sa�+�՞�4%���f�6K�������Ց��j1������D$,�+�>��H%��$��#����ٯ����6D���!��� ̼�*R�1���+�A�x�SD��%p�R���,8{&�|2��ێ�Q�Վ]u�����\�����m�"��.Mg�Vo�s�i[��`9�k&���tT%�B��F�f�n��R;_9������#'<Ǩ�B	����w�q����[0tE����<8����tH�/���r�Y�x�/����]�u�$9�
�ڴ43 C�	�#6i���O�g"9gg�|�ȸ_6����,�P�A�>i�)44P����.�a�����%�fP��)U�?ߝ�E��.Y��&��	Ȩ��E����7|�>S�\��o���t�S�VZ���o��q��?`��v�[k�������;��v�����+R4�+6߿	+[�d��	x��8��� �5��~A�y�7�������jёZ���'����t*��&�}Y.���nw�qk�p�Dm�����r�?����gH��?ٜ�'k���T����@��
:ް�˫�cwX����}�TC��Q�. 1&S��!��ii���u�إ*��֢7�9�?,�&Lf����,A��#�^����Y# G�Scbs f7w�X�0m�Ƌ��|�}u0NU������o^�T�$Fܧȷ48+��Jq�����l6�?2N6-8
�6��9j�WuVZ�d�3��Vf5��`��ݭ�38����V�V,����Zg;]E�ۚ�{
I�Ķ��<j
p��F��|����XE������QS�1a�0�Ơ�[�Mι��qv�L`�z��JA;����ZB��U��x>i�����CX�Q؇W�l:����lk��q���IQ�<�d��R�O�I(��R�9)���a���b�yK4�����O��a�"��n�ӎr
�������bU��|-*H�x]"�)N���)�f3�����	�^ ��z�1E
p�)j��ðO-����b�v�&�'COfG$dsg�E<}�nW�y���`�����6;J���B`!��R�}UE�l�f��+{jD9�Q�5�q���y�g���3@���c��>�1��U ê�V��m��-$pK��CWTI�6Rjf�(�#��w�@���aoE`�7K;v�ܞB.�"_t]i�>�n���{��-R}�A F5��G���Gx4��ޚY��4P� �@��� �<�MNT�[�@6���R]x E�Z��Nŧ6R�﴾Ed�LκB�8�Ө�\5�ޤ[\4Y�u��+��#I����Η�,G�g���.�N����;u����RK858�H�T����X?��EcN�=�q#�n+�G��zg� �#���/�;m�P��\�:�:�>��ߖ ��y�8��K�7��uki� �q�i�yt��;� ���:�	Lv����	���3aZ�|[����e��	�J��b�e~�������o>@�$�����}�S�F�G,(��)��E� v�vV��V��5�[��@mI���.Ŋb[J�OUXA�l��4's�aF��펞Xz塯8�#��(��-
pF#�W]�w���z�U�ۺ5��f�|!	>�_cD�����Z��[�+���D����Q���k"�%	��{`P�t��Tx&�0��u�G~������s,#e1� �I�$zC���J*�}�^�#���/F�5iR�W<�~)�O�2;Y��'����XJ9����t��#Z�q���=��B�"
=v|ܖ�I��K`ŦZ�E��y-����K���D�|r������_1;��@�f�e��x�AO����Ai�f��X��>��M�=O��{�=�ϐ�q�_ WQ�L���T���Pt)CRP��3���y�C��7������M�׌ђ3����	y���`UO&���Axbq'ܱ֯|=?#s��z6��7�3�ǔ�cF)� � �w�ޯfB�s���n ���ٗ_��&��x�.䀟�<'b,��#Ɖ�����rs��;�GR��Z�����s�25(�x��~��r	O��|����M6�Z���1Y1��*��RmԌ�q����1�b{�b<.�ZcZ� ��vOGvD�Dٳ��#Ă{q�bq]��=5��
��U���ښl�ךY�s�̪p��a�B���f� '�s����fu���Y�
�[~�����Y�Y^
�dA(X��°�] �������ޚ�'��5恴D���6߿<�Ld�d�)况n	On�_ŧ�헨虓����d���#�+��l*��A�s�����-]f�`)���gXv;Y8�ҧG�3��� �w`�ٴ�Ծv�z�(��Dz�SP�=݆ �6����6�&�k�H
���W�M�+
�]��nv=a�kb3����A���R[pO䤿�q{�aǳ5CA�����ݯf)�̴g>�G˵��Xg��~n"V_%"�`��$�K��a��W��}�4��@+�͢�h�O����Ū�|�kځ�5Giz�V��ˣR�ӕS1�	������j���U~�u�-�bJ*�~�T��k����@�2J�>K���I���\���d\=��*EV@���?vH|2�ȩ�1h�M�,:�d(�Vp���s����Ǻ�s������T�����:��J��������	�5��o����K7ᮗ,�T6�(%��D���#p��Wv�;���Y�CnG����ꏨ��L-�3O8g�o�h�w�AEE�p$ϱ�mf6�T1|��T�r�x9i�
ߠS�9[�J�F�}ٹ��ҫ�G&j���玀2ǿM[���������O*�꿰��ȵ��/鱔�wE�Dy�F�Z�(������,����F=<oWO�y��n����W@�&폼n:w�E����4�w����c�j=���"#C�SC�~�A�U����di��xn�u�/�}և�q'�������Kȋj{Ж��[��`�X6�!i��(���1����7K���U�Η���/��h��exy��?CQ� [��3M3�T�oI���	ލl���jE���4`��!�����5��Ӳ����)Wd�g����j�Z�3,�1>)��q�����a`t�DP �E���tJ��E@���Wq��YסgI=֮��B�F�	���; 5�����m�R�<�F'aB�H�i�U�]f��FNiZ�T�VL�X��^�Gw��B+�L�����Q��҂p�D��;W�OmCi��^S�>�qh�5n�Lc%�����	9��m�������>O�0��v� ͅX�f[x����ƻ��w�(��)�ƙ�8��h容+���+�J�!�����0%�n����5l7�:�u�y�r�3��Gy��g���!�k[&B��bit�Vl���[�N�o7ȅ�X�|�s���|��9)a-Z*���JQ�)� ��qx#�y`�|+�Y��$UHui�cSֈS`�Ȉ�a�\�|=Q��T1����l!�����^�].���_��ϡN^��ۦ�(�#:�����e-�&rP�%T��KG6=�9�!�v_����@m#߶E#:@%.ڄ!������l���>�������{�|��:,5:k1�M-�L۹!��>�|"rI��	��H y-qù@	(% ���!;��b*&�������j��Nztif�/L�M�ڡ%�3lv��l@t%�P�]kgc������V#�T���z�5P~��6h9�����dp^mc��5�Gc��s�߱cMq��� b����۳�������}��I�]��w�4�K��	U�I`Ez:�A��+D��4�,�*̊6�����P�T�k�ثb��h#*M>�)�D����`|S�r�i�Y� �j��Im�z��o��`���/�(v�h�D�
�|�?y*�C�*����\偹��{��O�u{���5I����Ӿ�  ˭�� �;X]��i]*��{S�J��eJ7�u����Lw;5�p#kI�e�>��?�E֩jӃf�y�.�7�ƨ�h(���%nP���L�~U��Q?���q��\��=L����s�Ը��v��˯s�Ɔ�����2J���1� Є	�뿣j|�I+��9�|p�*���:����M_��M����T�+����5D�TmM�'P�6b0�O���0�$c?;w