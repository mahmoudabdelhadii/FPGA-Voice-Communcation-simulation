-- (C) 2001-2016 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
R0RzcrNyKcl9kR+fgp6qKg4ofs5I4fBjr2R/Re7MN+Ut0iDorOm/W9xlBNrSdkq3AYOH4U10k8to
ULJpIe9RrA94+VALIyCXoJz1FhVi5VNIlqJrNmZu9EAUSpOjm7hQJQU7uB7Jg0wUyXNe81LKZh3s
0F5526W4tQJAhSG3NYvigCyHaKxk9IFWXP0lJSROGoQsg1ZTWwqcmAmRW+xI+oMoY9V/4F3HK0O9
0S62cqelGaFHCP0/5LyLQgqFOolsdCjZlovSeTfN0ICAXso3moY6Tn28E4GBx5CuyY3Sw3WTOpSU
DCH4JvBtOaf/iMNwJRsOC03bLHYlzsOyh0H4Mg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 24272)
`protect data_block
uBkYuTI8yCULzwqqSsLByPNA+AqyYYADlDp9S4yqiFQRCC9piV1/2tU5DEhKxX/wKdRu4KttphN3
tJ9YjP2afN5AHvhe5pyIJInej2EDIgY3FrEutwYFFlUrFgYRBKTRf9kHtyiCa3C0f41rUHTuCKDP
7HGjZ/doc6CYPBbV/krZu5qUt3jnCySl376SUjWasfwYUweTbwyBk7CzEyel+QMCp6ELgs1jDnsg
OGFhiwPaMlKo5d/HiTPnLpfY01g0f9hQrMBNyWNOVgXDzX5quDsCEA5hKaqlujQJ1CVv4/8ZUfhP
U0rqXmMOK2rbYkYppEFm09H3Ts6m++OS5L34MKkzd62OZPX6J/d3lLvLhNjXMyUmOqeA8A6Q7B1K
+QfLR3Zh6vL2vNB50NE07k2b1VtAx3klWYI28vKI+sLI35wVs3Lrv3odqVk5D4ihBkJtQeLQkCJl
1E9tRvlh7srE68meCBj/AiJo5wfnECXQrQnynVdzmvxKwW7lxWQANdF/4RlBAE3Yfop0blN8PrPb
4FXX+jhuK9+gjoFM1NNSI9VlXmSMGvo05MFpI92eWHWBFix7dLuUr/dUQJCqeaBnBBiSaNOjgd5J
5CaQvW8O9NZgKpVSHA6V4zZo+jPJhMQJ7+ai40EdM9fDXoYRn/XYqyGnIwjLSsuRxUPeWEIYW9cQ
HLSXtVnegipJ5RdiWXEyzFvwy5oJowyZTHG+GN1uY8Ku1dixh8PX0+u8uLWtudUrJkoP88kQMnKU
VD7VRVQIfTQSN+fJqUZn0mSGWHtvFrnohWLREqi7BP1l2qDZgApRXyx61haIJI9lse1yVSjGvs3m
xOp1dePavMPzfx6XY1hyJ2gecuOQhnegkx8mF+7egErGs8KOMogqzpFbQltvTS2bmF7NYhax1yEf
GWV6665H9GOiHgCwkeTopZDyjCxOPbWxtdaGcJGCFMIexXU8EYOgbL441n1kdAp/BdhlqHwG8f3G
oQKOqy9ve4sf/BIHr46OU32Yi5MrjEjtYvPUuwYG35wjFC6omNbw5U98sBoturxErmcqdDyTYMdB
hJi8V9hTzZ5hJm1/lsIw53cKYPt2jb+/McyKFSnvmcApcSE+b31lsdUJzci4r/pdLT7VwdiGZS9i
8aMc0EiAYw9n4CYmb1AGMmnzjvzGdr1GS+9kje0CAq4mPkdzSuB5n5GBdAtgeFA7dIjNYhLYABp3
vnxOUGq4MFZj4YdpcCjw5Sgtlam5TKBp8GF5vRpM2VRRk4goX4FKONbgEIP9i1RBeIVq1TtcoiSf
Pz/PgLvbSRea67lyWiECONeN2R141O3/iOzAMXOtGS01bUU5jnPSGLL19LJ6SZ5vCPKfHahY53tl
emE4ltsR2WNCb/I99ME0GT9lV1rmi7wmULxukjFLaE/DR7HK1b+RK3+i0O6TiC0pw/xaaWRwCpAG
akTHBPlTVuWwWhS5mrhrBIYEK+AlWyOJw0Y3Pez7opDufD6FNh9EsMg4RhjvGYy6xqrPl7JVtiV+
qRAS5W0Lsh27VNvVwHv5p2gSYGpETB9L6JWf3gliF2T1Ba6zOGXi1lY9Css99cMo9cWKkBl+dfCy
OixfKfhRDDEkFSs7r6Xga6V42jpttRCHACboHhIXk7xT25h3XqJe/W85dlmxGc75oZCaT5XQ6+GI
3t9sBDbchwK/X6oxCE2m9pK6ZXJqeGr7IJ0aHGtiw3QrUrCvzEFIEfgFrWMcL44Ge8+y+Z2Pa6+g
tbzlUmG+d1jzDeiVxas5MGFrra9HPAqq00qcAcMdpbObuFct7ZR6D2D+GbKbDRwOdkYfFErEsKZs
9nQA7z/tbT1E/b/T55VKLSOjfY36Zf08j7ixEHRJsUGIJS6ePwJBYlLEN+5TDPykcmik/P/gk0dF
RrgNB7ruq2912BmKcqVNVPDtlh8aA/B7FdMQwUPPqwvvMQbBjmJRq9cCfL8Me79wc0mi+6NsQDHf
37g2uehjaoModsmHaWN0/HikjKYP31PmjPeTu/QlgzXCcB/7Md6x59ZBMTtlfCOO3aYx7klvt/X2
oHkiyyqy9cJhzwUNQVJMGx9tIoMH0WiRus4omJDiXkQSrnhloIObO0/4Q5yLr/mbpJLrYmSdIGQB
JvFE/Q0FwL8osG9GC/JfKTlXKAlgf9Pze7xLBKQulIGLIXpFktFum22M/Nv7lwy9dTIkDMJVmT4C
jVP7HKBjNMo9S3oW2+6eSf0yWmqLH2kvvU28J1nBME/IQigo/HC/6nTz8ofLF+MAilciH/nod5BU
rOKE33qf2Dqlu93zo1SU9fwWZRX96vlRA142BulB0r1E5AzIndKY/u3B3uLINV2SYDr+Ej4b7YON
r45FJky4JbkwbnO0cd5h4sZIiqIR0svZ2ivw6U3PiJRw8SMD7plTxNEhE1gaa9LFRHRTwhif8Wie
tgj9MO/OTctolLamR/55yKjJaJWkQypAfRSrt3pGsULcqY5MNRAk5HdG0TlDlE7x/hTN0iGLfws2
y8dHaLi8AtJCnFu9GU3i+aGlE6R2kCrrrcDxKC04cNNtbt4JyLmEHHqDlrLHd6vLEHFBHt0V7zzk
PovaF4KLIuzfXxCYcIowx41y4W4Q2S24R3tYWcekG6pl6PguvqZ8roBeXUaXNpBYXyXrq8hWWR3Q
bFPtvlPctLhlkl6sptPxZFXaEZQwYiK6AyIuI6Fcx7/It1WyFKYbB302JDO2yp+zvsGurbJQ/+FQ
Nvggu4QKDA9wHZSDuDuQT1BUAWUulgqxwSVmHfMq++EuDjhq3jWEP/8fL4jke1+VsNGpVAsu6ybu
tHFJeGikYeiLH2HBggczbmLB0WvaF42hVxxc3bVQcMLPYKltCTP94EgMcB3jYMsjTEqNEmGs+z3R
EkyYXsd4A5P0u6uTCHwB5R1daqJmoVy5kpWD+3ABJ8cwnmXSRv1cxaliu4It+XHz4jMdKy7jE0d1
BTcKcPK7LPWJYXBFhDwSWhDu7oFfDy52ivotAAkAgKRfOcNFwylRWMmTdCFA5yFdtv0JSPugjwkf
qcsW1kAJjqUo6IHuk+PRuRAL+7y45Tey+M2zbzwYQXyq5MLiLzrHUqnPScDHGbGSZWjkomo7NfQF
h5CM2+JlyglsK7zPwQbZ7vwSNQPHVm07+3qmmzloQGcHCqPHSKJGOybWhirEOwnCcfEA0cjwFhOr
L9o3qn3AZUTQIwxHQtef0HgiapJLERugT1LRBsKqkbCsHtuysNcW2mVBAMw4zZWa03qHPl7siJE8
0cfK3XWRgiCgqu0nHlZ7BpFMTnuG/NGXCppNwMuFqXbJpZzmge6vXIehxYcBpuNniPwvooOc10m0
XPP+GW1mOSxOtcbvu0e3FXuju2qJ4Z2sHMvhTTcGLeQvntul2zfFGNTZvqdMqgLqZ2n7Ks4YO8dh
ibXOnrAjnhbnl8IjtbqHzlPKI7jZ+MA4+ZNDMJdYYzQu2TXo/KaBykn5mLmHOdbGdlq6iThmLYlj
upDrBQtg81c9Ob9WxmQ/cBYdNGqUCSyIY73t+ci8P5kwbSD86/x9EwvuHlN2Tyg8d41XXOmiqpEC
g1xmDGj+P7epiGOfdoh2sW3Qeo+yZNoVB3g35JodsZUtaZ688utwdb8Kgku3krBf/gNJlIBnrZWm
IuD7kO4Ts6G5csNWZdzzH/nqMCzNwY7OCK/khqtz8I5lXo3heC4mwZXjONE+28RchkdVucbw4hhG
phIqSYH4UEl+OeCgxXunbByLcs/BXdegXJNoQgXPkQzIKHUGQOJJ+kACyYnvehz8t5rF6O6bsqzi
2DSAiP/iLq4wnxAkaxK8AbWGpMCY/0eGtH9rOeKUH3NOGkeMjIBoMxOVwY44f6/A2WYWZJt43Ovh
lrlnzIpIT9pQR2zqZ78qynd2qCTUTTFpAaC/x9TeBVVJ4blLtBAc5ce/w3LFkhjKVmg5YIg+LywW
wCH2UcEn8T2qerzgPDcJrL8U8JEMXcTJe2QUxsROh1Y05zIvqNTFTIt6eBls36LkWEK5l7tSuKPp
TlUoeks7/2YkysCbd3zQBVs+VHNvCd3SPm/0AzIZAl84SPQE2qeBt7DUe9f806tsG048Zg/UHHpl
Oi1VW/yJdz82jiSYJapmJdktA9Xy6QwVTove5bo2qCke2lC9l7evNw/X0waqy+gy1P/RGTE1aIM5
ouk+vwZZDSh7mWqDtOY69gNeyeSW0U2znW75Hl5Cjcduckf2rrkNlblbZPN16E0Mg+otGqK9CMga
3uvvO9t9/2KIgKc9a60Rh3YAPUzhjaoRpVjsa9qpxBtqLcWcGGbafuY0URUOpEQWpXCC7p8Hiben
QvpFoJ9l01TNa0ddxVet3TDeDPQ4/Qh1hMVT9LDgwo3r2HTogQeQBiQ+B33S/Kud3RxqBguvvRp8
hbkBHomwdSuvD3a+tXPde0hKwBUy5awbDwK7SWDi3CwsW8btnW/VkyRxQfG1MzqgVeGvLNppVYtP
MOR8C+cMbIGNu7c6bzbAm24rIm+eyMkRzRta889BuFfPdbUhqQwNqXKDVtWbTTS3PfrfGgE0QP/Q
RiZq6dPEtCvmnqEeHyxCwCILlmGFZiYIFNh2fOVQFUJCZJwbtJN0FTf81vi9yhVDl5HIwnwZalxF
dmmoAURCXsWT1F/8e+EM0CJfCHJsu4PD3Yz+mwXgkgadRKuYXVbf5MEd4LXu4etKD6auiR5UkVKY
mFQwpXcdYsGtMRTLC2xdM8AwjlA6y6uNg/tD4Htaso+1OkvmHhVbvrZLyvwHpnYzH1VXa7VJmdfv
dijlDwy2E3EGcrP+nkM6r+fDrWW7FNWCd7lgo4aOae901kZcqbxrRh82XwtKUIzP8jK3i1htxZo2
MCLnTDqh2OTJwLrXewHoGv/VzMd0pylT7Q87FdjzdTaHxOkQdku8hq6HKJJcnWDJFc9seX3MaZTr
Y5cPTp6c7om1CoYdLM3Yz9q1y5I+32vgBh1C11c0n1LPo0hWOLkKji9lZhRKp99H3KRthlwJ/U4t
RqmB/q6YLraC0GdTsyO0qE+zpuTjOv5/1gelLNha23Scbra4iA06dmINr5j8JJATcofhJjeS7p2t
hMWkmM7r9IuA1Hn/m19FrvwCuf043+B7bbHhSTW3gIj0YMpiE4IKcboPvUm7iScvlnIr8HVXJRaY
c0bhvjrQc+Y58DIg3Wo9w0JAUMTQU+ZDm1ku91sOGNIbVcUDmIlS1AyvpKxKxcbA3Bp0/nDYaffJ
KHqYNfc8B0KvurJW43JxWMOktpOUNj1tZZvv9tjZ2B5pobzfsC1lCoF5GyAyyG4Ddz/8xRMJ1YT3
XnmiytDYhhapgV0aUSr3zDxH+lRYAJoX9rFqPfH9gsvZpysIzrEj/tpQCLDWR9AyDLqjsuGGK/5V
TiyPCi3gna+IgHozmy9gH5Ei3S00yJDKzR75D/E9204sbUzrllCnvEvjK0w5wV+w20JJkfG5JmGw
RsAtsethXZUkPhOipsCZ6JuevZpNOSMjhcPmVHqmIbW62V4lwrnQmjqjQdmnsXbD1mudA3+yBRhz
Rn6oFGORgh9GuVeqFW8klLi1/YgDakApsCll7+TaD5T7D/1hToovRdEcIDMpPbLfdf5RJiTbxOca
ZJDnHsVyygTkPLSkwP8o9Iy9JQ+7nXT+N2bOJqEDsgtgzOPyRVR82a44cphrJO5t24qKO2PScvMc
+AlpXfoPxp5yrp6lcYVcqkBI606Lf/KUKW08nz+HeHxlzLadsxZg6Pe11ld7/njEar2GKAite873
zUEONs+f+ef48gOErGdEV9uiN/rIeSgksY+tD8n01+Ua5TgA0YxV7SLBlQNLEgE0uein1BG1nxcP
iw/2Dlo+6Nv8JliZJ+F8ejh/2sfHXxG1P+FFIj9jYaGpWPzE0wq2ZghC4amCK3wckk3z/kUKqnlt
vqGwpebj16yYlPQrWk4LvJwu9pZqYsjCXgKnFUihrj/XLifat9yBUqPrilCqexoSqMjOR1T69EJp
49NcH6zCkASs06VmB/XjnJGTn2d9f7IpeGUd0zcoWzifw/MGOrGr7yBHDP4o1H5ZSpIWwvkuzCu0
uHSKgf7WadInczFQj4+7LNLBe69xWqCAuTWCKhMn36iP4mBu2H7Go7qcTBRw7dNdRnPWMhgZs72H
hSoHbaN05i0JHWCT9vedpM+F1/oOR+IrCnsNYVFT0lNt+p1fKuNl9YX/RbL4yDZFg6eRrx4Gy1ab
Yv6+mzf+XOSFW2b32EyVJeLBHF+D8l7ut5sx8zvPT7WYx05frkVn6Mf8gBnplnmRZrW9/ppmVmGG
KKyNJ0yn6YWs9hCp12U23PV4OUubkCJtgrWUFn521x68iY6ze3Kwt3KuwahW+QErdCJ1bNuQ456h
jsJG4yEEgDZy1IvBf1J2ggwnI4FPO0T1w80jbYPuMS8WafpbA/4We2/wWrF7Ki06+5fDLycDiSpa
xy3yGNd3Jfn5Ah5PEImTbdYsgpzpOrQ+ycaB3ZEe474pfRujLf3YxzamLYojN7dhG5/RH6XYV6YZ
UWUaF4ptj+xtgkQ03fshmcohRYh39CyPfnKVex9RJgKhTuLl0h2UwijMvuCSnZXEPRv5q0LT4OxC
dD0qDUWFDsDL46ZaOZvRoMWkIV3McC8pbLFBRZkCwKLXb1iNsB5c8M7RrIrgh1l0df5hETfQzZ7J
BIjNqI0VxH08o0KBvpeCd1ZFGMpmW/8Q/R48DRcpRYesr/MGgnDfhGA8dJOcM74IO8GQhzc7GlXO
2LyalsrPHRO7xKYznFMHztcG6TuHxLLNbQ2l5sgOonSXG6Lf0eG2ocg1crOLS1nnrSwTVzgz/QO0
BmlKTiSjfzsQuYryJPHwz2dw6oXzeTIHe8QdS3epws0sDQIbltI2x0G9QKaNFnbUrQAH8yOek+NA
cpOoFzKnkr+7HUAINafpDHZXS1WGGkozEe+w1RmrCW9wUDErpd+6bibVR59dhxSHK3N+X7Rj2A4f
A5LcUzFRnnWYwaD6v0mLm8u0/emNCoDc2ACnfP/FXYJaa3GzPdozYpiEdUCivbdlOGurA+rFyQRv
u7Przl0KkVwYnjsMVVCqbDG6CljSuIW9QWpXMrW/BdaIAhzbJ95V4yDcjWWpIg6KYRCkgtQ0U6Pc
d6MoeuV9CXuafvy/6aizES5hL3AMGq+s4pVGGMkDOC8ZUMjm//UpL+936CeDoyh+ndmdLY5cSzwp
VV2br+CY806lgJ73u/PToVkJKhzUEuDJyjvM/acNbk/HCXciXQn3YuksTEZn7AFsvDgnGD4dK5qU
khwPH6M+kwj1Bb037RL7Mj6NF1imzXC9Q/93HJMSRDOygD4+8c0TDfBzCdGg7VL5cIheT84NNDnN
/jcuzidXVRdWc+aSxmBsrOiqYp6xShTIQE08m8RL5a2NSqnpv/FUjbKpuJOEmQaNWUoC1R154Mlm
lVBntq+dRClPGb0aJEA3iwu+2cob2hXp+KmbXaVyepYi2dVyEV1c9ZYTRNlCnDYxl+DCecIFQ/4X
JlhTpB0IcOQDx3KX4zSBtKXJJDaA0mePiB+axEB7d2hewbkkmL9OXjVXVcu/a7eo2pcH6xo8C6IT
pbAxbv6CEW/Pq44lK+prJwHz+RQBe5lo8K+Va50j3VVZiixJAsh5BCWoVapPv9xuEwELnJSJrOUt
nEHh1pf0BjimPuwgDcDU6oU/4KR3R5hyi8t1RTr4MH6fN0wq9NysItyr+wbMLWBiZcaUy4KiwZQn
T72pOdm9ntZ6KN552QdruZzxg9hQG/RIAIcRav8qaKLWYEaVTjvQLt6Yrmfe39X/8AQF9WrFzkOZ
4uoVOk2h2YsaTkdvY1FIU4NywuuYpWkXej4np0SL3mUQLxEryYyuWkeOpV0v8FMMxORQptBf6C7t
LBVRnOrwCu0OT2Wmm3q2tI/hu9WKaHfDy5QvM2qGDqlsyOiNU5RIcoUb1Q29fjzEymBpn0ywE84w
qyyeBnCJN+t6iyuJ2K7Ksnk5p4Wjyej/F/Q6Hljd5w6P1KjIxSw7GhNq1UF8laMjY0Qu0FbM8YUm
yS0X4nJr14OajZabovBhpY7MOB4wAcfgWy3M0puHXKgBZ/FkTsHphv3ToQM/JAP57Lmnk9WOiR87
KJYbgyBxu6jvdFEYYTP+HAHTF8erOGkwfIcVXAVO4XY0VndHbG7NtRsgeq1VD/h+4tuwlNDMpLBJ
rcGOyh/E3pq9sOJJQ567e8uyahJR7G/R92ApIYbCbgVWDv6iwgtlmXV6YTp5aCWG+PRbJm2TYAr6
3Jo2m8CV53+9ZpOMGdzuqI2ZpmAZhGaeIUOXnmWrYLF8BXbJi8P8dc6QE1zTrJB0fwQ11GRY25Lx
Nk0F7mW7cNiAaE1SjPCtMlCUmzyIpQMonoo9FwDIQsf/5eESkGJypo6ewdbZuO+3ncD9V/7fRMIq
pCorkGU9R3HMbExfxlY9DGZeQcm6hcSpVQxn9nMeDF0qHA7ycvDsQT6NVdFdgdAa28HOV3XdmFo/
pR8De+gHrmtktVgoAvUmaDpgEzNqgqJWbMCYzrDDlad4uLzKNgMWVx8nz11xa35x2e+lHKVQrn2V
U1x2GI/ck5gswlUecxVYbY0idgDh+BgdYKTDIR7q0Mxu6evoFjNZsLz5lPo/B+TxzJGORSikD+Nu
VAgyUzaXqz4O4SqLwMthbMLMkR9S/vzWc4f0+jjUUGm/KQ9YiqluAN9FXmj/RHFBYKFstzgoSbDk
St1WIko2eX/bvhZJWXeKTGGM/uhLW/7YomQnZfuR/KlkXq2DF0/yyIv55nTthlkSecqwWTLYPxVT
4cjZ3WsGDfwmNE54pW6gQ2vMqWJaxD+6TUOg8kGrwpUvms8oZ8d9jU2CpXzhDhXaA/7aMudI8qCT
+Tsxek3ZO4D77C8/QVsxJeg3sXueAhgfdk0Ozx1KXWuw+gQuXYSA/xC4uK2U5VsBrXycUkFjia2z
+NvxXa1FBIePQFhLqGbYCbmihdolsfBBV3x8HGM8PVg/jwSid7YMmU3rK//Sd+4zdObyntr24KoI
wK3h6zR3VJWum1PL9z3osXsffjXWJOskA/9GOnEPTD97rq0HEW+jg57DJFBj4OGpdlhuZsIUEJsB
QdclO2smJ7ECqGJLvWml6FfwbV+8YimfCjhWKqEKpnsaKLtJYPDzQ47h7lHFNfCrf1082lIgiHHD
r1x2YzDJvz3rxe4EnGW1I1weTa0TA/QPc3YK/hHDBC3krR3rlr2N5Wj1AHA+OIuh13OjaCIPuO+1
OiurFSPc/DPgCDQNpnneCOkbHfNF3v3n8HU1SPi6NP9XbY43izpnwudD4QsZvvLHWsCwxN7KjQle
Mhtx8vMgf2KMrqkNdNHMK4uoR69ovJPlkDoTa9lsQnCuvhlwdxqsTj348hhzEv7VgSgTOURPZvK+
7Z0i+vGV+gmbRYuDJatGYVTHgTvNdficqt+nYNLO7G3vpQkL1lR3bhyMgCMteECH58DLQyv6u/RO
s047OcgaeLnZMkvEubQrmu0LOLJc30HTHS3KFwQpXfJjCmDmj9B//5o7ToI2TRc9yD5vLqlVEnsi
dISgXbsapteZGIvaoU6SrE0yxLX05GkxK6wiRfpW7k3MQ3bOulyOCTDkujvPGFtJR4zK19uG9Z3S
Fpqr0ODmG8bUXGqwRH34VRr8ZUssu3W8QEr1zSJs/MjDR1GFc/FQIcawd/1JLskZoe4Kuxtkc6HF
e8/cnq4bLmJLD9+QYuPLzLAOQELI/gJHpx/vlwCxLFmo0TYOsHDiyJnf/q4sd8maR1U1kBvU/t3r
y9CZ1GaKMO10z0KE19jvf5tkpdiQidZ3acRDMLJxCneQeHeswBmDEIvfeYfoV0oPx5GJsMNneTkt
In4g/J470wGMa3R6L0tRPjCj4TOd7YdEjXj3bU1SMBQwMgCnTwALVtlZf2MP/TQCtiA64z7j1PG2
PXzvDDd9RTXqmVBXLLndfmElx8GjAJA2468vV2IAX48+n6b19s1bb1s7R+QXiqyYBbIte/lvLwRt
ra7qGMGZA2PED50R6pCtiM5laeua3ZF9pO0NDEsinfItblGcsRAantFT6X7g1yiQY+i9jhQ4CzeW
JfnGmyPt6fhJfoF7lUgzMyZKNyhtC7qaOby7lFzClgQN5UUnT6uliNeKYGUt/eQnYYuPgWANpBA0
jnA4T1fOhMgoWQ0FMJJMbywmbwFtLKXJYADilhJYGvevxti/WGdnIqDKikNiu6FVgmXl2+rZhakp
eQDIVHbHDp/MoulLnR+8oLst0yek7/ESejCenq1ZPvGEL5Rplw9nWpgEyB5fmPkWm3te3hvvH5MD
PyDmJlCqGsV2PD9z0OEOoTd/6tG5j44rQA14AFRTL285+2boh9xG936v/flLA8izaRczPAckLDYh
lCs4jP0J51+6a50pLY/+4bqnOg8R9XGmx2d9ypraLqFgnO82ZChaMBl4mouPZfdJzNQ/iNPKIadL
VrN+NVw5HFQIsj2Zlin7oaJ7QRkrSa/o1eq+KHYMwN9WkUPpgztU/Gz3xFtS7QoDWPU9sWGg7LeL
FuMyQfay0tBbj2f/zxc8akkqYJtP3UoVTYVGj9YY2s0KNo/H+gtkolObJ4BdBl+h66tcLS1IlEYD
FhayiQxC1ly2KWdv1FWc6DMSsoDrVA9eUzDWM6SLkiSOfzmHK6oy8W3EoIrOYh5DNf0vmsmVC1pJ
LODa8kfx1j2xzqJw/4357CGL9Q1dFsZoYFOQH2fL0kr99A71u6vDu4BpLlVR6hdhxbTbwlA1g5ot
/m5G3aRGQdb71Fx4jLGH/Ou0fikHb7N7nMpoxyqhfytHw0CVZ6OmGvk+/CI+IhAVQ16iMrviHnAO
cwKQ5mH3lxJaQzbBco0PVC1gI66KmtrOk7yxfyDs00jDaX5XPEWazOGntNmWKxbnOsV97taDl8V2
hrOT4oe6u5Gu1bHi2mlykrg1hzI55viJ6GeJfkYyP4TXqnx3mNrvCcNVDesJeJ+J5YEpcjQZ3bve
We0xdLA1pKDH5zCyr47i4X5xufmK8GkND4dzkU9vJSmAhlJ2SA+Q5pz2wYrfZJFFoP0Fx4Xm0rG2
Uo886wE577JBr026ABLALfwtj0hVe1/IJDobKm4Q+AmH79f7VkdrwOji9Poi0+2rWNjy4oxUliJm
SqQRTAPix89YQj6g4CcA4SHZKEpashad4ZdHgDbVRRka56bRsu038WEhv2t2SEqWJxcpteUy3Hj+
8r4c1WcPNJ/9Be3fQvzfo+xHK9krF3eJymEUSpXfCeqGdAq3PDzz4E1+USqktcs4/auWdNezudq7
HyDOSkYNhsGu12Z4IUFhTJM0oj9EUeK3oX/x/idMjdasfD8FEYIsKrhgrvZQx8LWrQq0hR/K4G05
XZr5dDJYkvDuw5p6Qep4V1Lpz6MvH1h7dqsIH5wBs2+R7SXbQ7WJKIlGgbO+wOaT9A+ja0d6WsJJ
YTfgBOzR5NzQ0i2IB2XC5SxA9abi+wKyzDw8i1PFrXcYjbOH2o42ozP2FRI8KYKqEUNYVYz6dxSU
LERaEfSIvivxslm1ZzThdrMdU5AB/xYYQIpMzFb+WzfA7PaNl8wZwwbxkBoGr7EqTGbS1ImyV20e
O72Vj5t+D0HeEo5RsFBqIyh8k1AjDab8ANx+HGmaZlFyPOgLdlC66l1eWxj8aJ7HDMy0UX6HsAeT
MwoX4kUKocJ8PekqskWpbHf98ysUwsjf0cQhaaPTECyb4KnnneP+ERNt70GEiJvN+vK9BpCFaL5M
pbab3/T+4RaBeBcVFKpXE1KTCfWUz6ts64XxNCcFSkMkiO2oTm7Z0TqOle1WaJgrtZbYYWViZWuG
EBQPp1yn014Ppx+RyMhg9fQbzTQeQbHgBfLxfg/oxbJZG7UFSAn1gvj7eMlm/fyi1m/V4ZtPJxQh
zy2HSjaBiufbrueW5hSxcEhYkeRd+3jRp+DsUHy/aYjMV2o7Ethz4pi0yuxrv78mz5rQgFs1l64M
JyctDrlzy0x5sDTIi1CeFKjDA+Rt05owkhnAIMLstVYYsVLGG1Hmed5H1On+8z5liAHfCcbFE/z5
qQs2kC8+ZUM9RCw1GqYm8FIYZd2lJKgx5nwjk8USAQDqksa4Fh8mn2hNoD1I+FAUeadlo54logzp
ED3y0nxTRg7oUItQ2lUX3MbR+tZaOyZS/S5N6dV1rAHLuizF6PJYbJEuj1am45kJpnwulvlHPAnP
kod1jmJNQM8n2d4rAVRB3Vsav+sVhATOHdD7t09QvUM30+4Hz9mtunkg9RwJIYEliyzTVXBHUFHj
4ky4zg7HpPoRB0suMtYD0zUM9bYql0x1pjKRVh3/M74eOwM+IRe08eJD6JMMA6xegvhtDYSJueKL
r/cjOqlHISUnAnmomt3TmIe98iR9gnl88mGqkVaJOsA8XrConTlQ7DdDsSAvvC8IFa9MIq4WjqLa
72KCdevEBcbIgI8KoBWPm02+CK5VO+lAiQaeGG8t0TwMrre5VpgiknoaRPct64zhVvVuMA+PshbW
oHQhNNK+Xf/73Cpqzc9XINZ1kmKrocy/zI/c4461D4tiKTvVPFjM38Ol8Kf38nMqHc1f8WWFD7CX
D9z83+acwz/CiWP7Zb7EF0gKo5tlDnYc6XQZO73CkwhKSywb+E9Qg2xDuZp8lrxHjrJ1OzPxQv1u
WbvpA6+dd3f6NhUxgu5ySdD1/qbMUSdZzPfcnPKSfBoCa7h4fG16CPUVJW+iyQMkp8c/OATYAPnJ
5bB+vUJNlI6siIwVPwpqV6hCeA5/1c52gV7ceWXuFQVui/1BGd4x3umnRJQlkFiKCBlmYBW4Vs8w
wAw5SLeLO0GVFqA73S/txFogjq3826NW3ONn4uwWoOR/Dl7ZENCP8lFRWmaP28tEDvTybDQtkjGF
peFj+A+pBHvVpf6g4S6ZYaeqoyN7D2r2mWruML0VYECrnBIIaUBenF/w3Qnw1TqP5PBOstTfGsfR
YDOI8uJIs9Dq4CWRs6NIp8GgYVpT5Goch5bQTYiK0Y7mYIQ8ddU0+EXtDrpLVhvWsUK+johQEze1
MYXQJHQSIau5GGCqzaL6YKraE1jSfRjDZ5QTNMkZT/AlUoMk6NYx+etQciiVWEHfGqApVznNqwD1
MZF9dK/UARcZNdBrUKY9PBi+Rcukwqm7JUu3ePFz+6mIvmV/GI6KFIyjTNtiovywQhbfhiut57Cu
HwSn1mhfO0L3tSKVP+nz9ZX0uc1rMRb2w/wAa3Mcam9fYuOOv2qYkrC4+rFVEAChQTcM+COVo1dn
cFnclwq4Df2g/DoxDloNpNYjlznJfFWwSZ9M3NsFdQbkQN4b5tBxyjw8Cal1dt+htQFjY33XIKly
NrKvcxZOXhGWSH5EivecE0p8D8jKndimr/E2ZPTa3Hq18WmRC2mCEQ876pfAwnmIH7ZVUQTId3EW
9FOCyCqjOFR32mobucMli/9g+Dz8WC79/WczdiyjZOyD4AQg5EkpnOQvAQbvvYwRd8Y/ydoWvgqj
L2ZlPZqWD80wrARyatMSjriokU2ZANYsTgZNQoJE66jS8MGyfPK5L0rY7ORs2KmyGX6n7htuTlFV
Tg78nRNu2QdZNb9dxal289QvWLCzdEuE4g7oN3dNwupHVtj6Mtum/y2KRFudjAtzlUVvj8E3bf2i
dmFKVITgjY9A1YJzo0pT6CYKH0f1BhI0/SeGIGn56or7UfbiEg8w8Nb5NtT65lVx95St9WniqNfT
rACqzVk8K/kdWASmObrOupy0ziXKFPsG7TWPRdCH6niI4xUp3w1gJTiCVqFZVpOmwSMKrNwbNfyc
W45biX1WspZB5cwE9k/N8/5iBLV/C9BMdu4Jgzpyw8E5RrMoyAOpqb1eoN7naRpfck302DrJA3Ga
nGxRaDbWeNZ4F8U9KYWRJX7vZ0FRIf7AmuX83UG/IUwK3cbOPgaYfzu0QPFDwKw/2w49VC8emlqZ
uYZBcgaDpxnyjc7mmhDHmDFo33ra54aPYXXdE3KShqVkEWGq3DpmvIC6xmBJI2U2LmQd1Neypt0k
8ImACHen8G2/tYyYtmVGwVWoeE97Nof5z3HjI7ELdP9wZW0JTxp+y69wzaNeHlroeXGoU/bef6My
lz05KliwJ65TpgNyxQy4VHb2XtHwdOSSBm7Z+0ss0RWzJrZnsWotXmaYx6hUVDuIpRCzspXxjT6A
nl8LSxTXxMQNY5bg5dMMHXSiI8OjWIZwILyCm5bFlbq/JfeqzOqPe6zeQAlF2wk3hf7VDxbFc62v
N9QF1mIAHDXBeR+JQv4W4Gci4ml9Rgf8KA1VSft0puSIDOtnglkp1/8LzUhgW8hKomdd8Oue3jqC
XyrIhkCGpI4/DLC66a0QgCC8SWSendwpznnYGlx4BHfoRpXz92/ukvVFT1dc4r7+CE9uoGMbVQDr
BpsmxTP4z+FwBAKl/XQUMR3P/SDbrFvcbOGxZKe3Lll8Z518Mtgf/BYihBAmBtOQ1EDuoZKbb06C
SyQ8wpt1lKWN4C038Zz6PVaqTHbgx9ay+zQeqss+0bXAoLjQ7FTkGX2YGHMAtGQIWbZK6E3r7v0y
yZR+lrmglP0Dgz24MHvUPDyuxw6/+FGQiRiwyjzodJcEs+5+0GKsOpYrrxW0cchdys4dqt9zU6SR
osJMfIX62w56Ejo5votUfIXsimz8JcUOLTfJ5VC/ypXkXmqqIR55qnbC/Ks6o48GHI3PdsA/MQxI
HcYrbPHhET8+9oY6LfLY9F2BKPkGXxqabIuvHWNHDCt4B7FGkWqqFr2/XcNO+qvpfxnkT6uR6MFd
GPs6X7pacYdGqzUJdzJDPeLwe2LgDbbKV0EpzG/YQArhUTkAc5Y+jh3qvZKJAMPSvZREPtlIWeSb
PKWmte3BDXwMMpg+wv3puvfZT1CKh1b5HNQAwARFCMwIWObwLRTy3vUs6F6zrPc5VyWV2T+ZJfs0
qbH/m4TLhZ/JkDSyIzzFF6G9lAkNSGwv0bDTuFwf5VnaYDyomjQjvD66SiPeKNsKfOON4iWbh1BE
tweGLciooVmIgEEwyAVHSnZHEPUzmQt1rcmY4P7iaJJ/9J7wB4z4aX9DRHDYXmb2fQomJN1wx4Go
89McQONcjSZ1zGpUQ+5ny5AQB62iDOPJuV396ySOuo2EW5ApfnWguktaEpi5HHVRMe/NZfFnTpH3
r2O2TGXj7OfiDj3MIfHUKKKKTvEDITiaob32yixzayMhE2SFAuT3cIgzQrauU4G0ZH4GO91ssOiY
7d9EAi5NjfkFGwe6R38r0mItXLOleEUgrrwtSKsjJ6115pck3yCBQ/VQqe1pzYTWVCQJSZneCjr+
ZY5ulXqDqpnvizJJ8HeM7TJkmYBhOVBmzWdxi2LF1+sxnKfWUwMoLQoCvEOFLfWYn8NiU5pCw/GD
qpXFF8Frgqdgmxh/mDsbdSUZCSnSEJXuwLsKXTRPFOnf0dY3d2sc3YZDoRQJjIpqcfbIY3yLHQyu
tQsJGMe8+VDv2rVF5rTLd6eCX2TouNVTFrTfeXUjYNdfQB3aTWTnOI1N3hpzkKkGltP9KAnAUCGP
43hFm0PChaaHU95BitXJVgMWULByFXvPswZ78qsK6+e769ej96tTFAea5wS4Vs6kBNUoyhP8Fc2p
cYnvanWPfkAJaErYXwdpGEGYJ/1nNt39sRjc3LMI1e5xBUOOfIN74vxgegValOBGRtOWCm8r1sRM
8pzcifdtfq/CtUFAKAkcgllUf0iVAoKxh9MfkgPVJHbkZtQPNhCVCjIHsR6WWnc3SvNpJ1a78r0P
raB7O/rYE/wAttEk66FNy41+CPjV7gRV0/kRc6++DwA/gmPD7oz4zx0BiplvI1V1zCBZJ4EnjCP8
G2jrrDrR9GQuEAn72P4X9RIkMB9X84YHi4mT2etAtQx3W1JBFA1JjfHmXBlyvxMbJeDlU0gzAHdy
RFBamyu4CLZO2pte6lSlwMPOAgSYxMra8nZS2BOu3Ma5WGvd3hCMW0J+Rw5zRQD7bcb1ULSmUbzQ
Rr7qChDFOvOd/uKj6ianDlbuTBW67djwFWyYljMD0JoZYI+Ua8/NlqdJ7hWpebKbMsQE0yTMiCRq
p9rBEkrK0ForcRy18qoF7faj67bP0rD+dYo1wa4z+ORvpWV6PVcijsxTg3cE2o1yJg5zI2YQxals
qswW7wuZ0tD28WAHHHKQMMTEIJAc+BAITFzLMdrvwLrQgRKJmViBnSohip1YQ6Edgo5ETMeb7Moo
qQmeqlAHqY72ZnszGWozMFjkw5Tn3UMMQWqpqrm/tI6206bVfXPrp9PTlF3B8T9Y/8R3o+HetJAI
Nx/Ualn4ddBRnU/0/5fUXs3Nh4N9B2m88the4vFPjFS6PpQtz9pjkt50xb2OW/jL7/HHbcE/N5bj
julu4/5jotVRnabeKffXoXoeFMhUWXxPd+HBpTzLkuk7P4L0we9FWOxhxSykWx/b3ZIBUz07kMBh
5jr4w3zkq6slh+uc+lp4car4fw3fXyzZqfDhIeYnMdMMYUeWd24HhrbRav6TUIzqytbXREz73M0A
6u77/IwQ96WONEbLEQa3M1ncykcQuQwacPqlmujsTcSiSNahcOPr13+unry6QBw9hntHMiQ3PQeu
YrSgk369Zls6xx13yisN0XsZMhPJKXSu9mp5eBq346R9SW/9N2Sokn67CxsaZdFU8xNP+2NsMO3w
XXVbnV5m0SQJnbgpQLOenGDX3+oH92LovbikwHkdLJdM6ol+R+N4CtUJhfB6ixNry83PNlqUrLQr
aGRKIAc7uZHqfilMXAwwg5OF3SAEozNsLWYTD3lgf0TfmCD1NxeiUe9/a3gLio/Uj5aVRB8Wwh0J
Jow1lVJBTdsmEtxXA6NpTXaeXrZtrdJGMbOj26oNGD67mrn6jQaqC4JRtkzSA3zuXlyLtKmj8Mtp
sW68TjNkls86APg4wWGXySWVGB6a1SxvOtAQxQVbc+932gVwWQ3zfm/N4CtDdMythXE1UgljczNC
gVXEmkdjUaUkmMjojQzNt4G/+q20YLRHdftB4Az/Q4nu2BqemMgh8jOen6hsjguaZlkocJ3gxSFs
MVuOY70Fz2cdB19sanSnEOwuJ/wIeI87yUn22k3iKZGtxxxAA2oyEUn3eaTBS5KECTN8Y2Lb9Kur
RYcmieQ2urgpssQ/6Zvks4tEGBKQ+5Ui6z7H3sj1bN7FaCEKPey9BKUQIn0l+UbupKsZw4TjovSV
gwMTuQvoHW1hP911IzVp1DWrguFta60Fi2Up0mERrpPndbVpqg4c97AX82MRl8n9a2cvuZCwymUc
+u897knhvmr/gbVupQx68Sk4mxu0PoY9g02m3pZJs1y1IitfgNdC5YBC0Jd0KdxlOYASjLUzdvvZ
7sa9ao2bT+JCwG6qNdae50M5O/R5JgDnTL7u+hZFtsqmk+1tu+wCak1prup8Cui6xbzcYO9n+g35
6aVrcVNX+xv0pfc3YZVzk6+6gBJ8/HNCtW9x6yYElSePhLwohC/rZGaNQkl7Hj8GtlmfaOsmBDf5
IEPbsEaopkLgFUvLf7x/5hB21CPwuqLX4fnQvhASDMXPVmevjVfKaBqytrXAumXUrM06wbGaYt+S
gQ+muDtVvQQe141yfV9Pr0Z0cF3ws3nzvayXVHd53q1t2ajkvLU9TiW79jwfcG5RBRhkH5abyO89
uf8ELxkcplEyQJlmZTJ2HWpMRW0HGTQoQ1hrShwCxLtsj9NN0PaJ7AuBF27yiysLVApH0UDjUXjp
VQhPpuoy0E8VIdYCfrzLOScTupIAasvHVJjOlmeX0v7cus87UEB5tSV1vpbB7hElWbZ+n32mSydE
jr/UzI5rJCM8/K4yzemB/uoIv9WS57EidI2hifuy9J8Ri/WlY3L7oSev08+SGbCebJxBIOgBrSb9
yrlbsxmlfpRBfCp6aE6tZY6QlgQuBm/zq/1pV/KA8mlzdH4zeUVvhhaDdCcUAWcSk0bC1AZD3ut5
nWM+WUyic/BvDe6LP2FPmiyGNOp9aTUmXBji96cGyPC7jgeArHwGpByKZsbrW/o4Hv0p/9VhE4wu
wk5YOOTdi3NZkvoQkqqbC16thMYBPFnec+VEzVktpRA7BIjOtsVXyKwwf070df9xlY6J8yJV0hgB
aZWxObJDa4Dd4jMfzGAzqVmdhAht0sq4qOD/KB7qN+E4kwUVMfFqR2qCVS5awte+r0O7aOkFN7Ea
lCCkJSHbPYpjQy+GzgENg3D324V/w2+/k2WX0gTmFRFP+OoOfLXDl12wV9xrfH1O0CR0cfGvfjuL
gyQmsBYdwEkD4g38geHfvTCy/+FL4+0Y3mbE3nqDo5Y3fR7jjrfVeKj5/8nh6fbDCWnAslohZ22E
jTHwP5lVIoND3cb4vvmUihqohQ2XyBSIdFVAhLQaepdouGpwh5LzXt3RYOBYzPFrxXpTVmtV0z/D
ALLGOCCw1zjdmMPjZVIYBIHhekAug74vC98dRU0OVctYUmL4P7Cn2cvASR1Q98ei4T9lqnOE0gpu
c2mT3WqhwTOQk0cKWncLBxN/fpl84TIWoBeXJwYiZjpGZZoRQL4S7ULCATpiYMA6i/SkvcPIzu53
hOxzj9wMyPiE/aeMv7iK5blhFHWjQKyJ6PNUARDM+fEjHAsEmapiKBiss8RvVmeD/ifM009cx9GI
s5QZYz1ul+0i1MIa0eWiGJ/zGxu8uB+zjMoYnY/a1OWWnK11T5I5uCbm6T2s6qvpZZkrxWlcYPhq
6IP8ac442xzgo9g39iWF2JLIkmBofrdpDF0um4ojoapfZjPRejNj9+zL2jRsdhI2qf2vNqo09O8e
mmwPEjVWSXN+2a7j3uNwhbHyM6Qi6plYot7IGkehCUrFbnKm/wZ5wxOHVgk9dpGgODgaOAYonuoi
VvKc+MnPXLuTM8N3scb51tzGMab5kQXmQRFa7cDZZcHST2wguIlHaIiL7c5wUCm6WtkV9RHLSyOB
NcUOZG4k4Hy8H0gHEtaZyjp1/MAUjbym4YbOxlufNzRiyl7gWsrohkHtHd0/yA+JBLJ5kqO9S4Ni
VpFTLkH4f05x8f7kVNZbmDPFIg/AVJQw7UwSqxzFwi1YQ5BB6+FDF0KZ51TL4gppgkbXs+rZPFye
fOnvX0haUbTJGT4T2cEUHt1TxSpjsCWyxASnINWxongn+qZR5ATN2Sh713+RBSRAurjy3xvEjXfS
JGRHBzfQ8SYcEfNieeTgIyKHU9C7sfOWeXKsjfTbQ4h3ZhuMAxSBq4vFBQDMGfkOQF4398RQikc6
1zxJ7O7Rwu4qRVyUpRM9Yp/otWsBAAsp3bVdyTQYJSnCpqoGadttvl4WGNFpP13GEnJr9Um05hnw
iX0Dvko7Anjwjl7TsBm7fqSD5UTzb3cbT25mnjb3eNe9+QeyXdDooKWx9wdwFFb7zlN+z/LgEXgT
/qc+euk7IIXvh+xlW9jW9aKv5AnwbX2r8Fxpdnroi8dQE6m0zaENekKGmu0IUcZEagcWDBVlZHC0
KO7pZrv+8/fD4cUz8X3tOpEXh5tctavuFkHLCRcuLvGUFnWfB0+jfuJWBs9Osz8ByQaprp6++sfV
wRny6AFibruet5U3oR3O45V+lNpON95B85NKL6XmoITgJ6rpLk6qTi7VYr+oIqVGziOFQGK1+FOF
tGtWJ62krHBEiooUCF0PcRnYiuUOblA2595mgSEc4KiFVxwaukm0s7CLJoWozdsWBrrPRvwcr6yT
uX0bALHziV2fiwDajWTsZUvZi+fJ4wZMWDzMuLoPCSR3GW2h+fKOw5HvOe/0GcNyLSdXFMK9D5Je
i/sI7FQYQemBs/KMisW/xdTlZu+NBlXWHyLuFnLHvA17LXDSVouGohzGlVHL3c9aZBg3bnzEH61L
QO6AS2bVUWutodwct4jLXSBt7Kx3CSf9FzU17VF/qsn4mu5s77CL5S2uVC8NTArkumdlZq9wqmOT
AGTw4f5d/sZ/NfQph0LY5sr3q+6qz3bg5XkTnNcLbSr9p7t5IT7Q+T0UUTTXb9PfgHOcq5J8J1xc
utrbfxtzMP2/oTOuqrlZT9uWuwuvhlspjrzIKFHwd/BH/h/AssUzlVcDG0d/NVov+zTZtnfPFie5
7SkJbvY3hlvosIWdWqALF9b3IEmru/u6itxFCz3SOG9AHsumG6fmlNmzdjA6ez6cevJxbCxyfu1w
vfBtBFY2hLWOUuxapDNiqG8wpUQW7OjQjQ5qcZ93dLqTZ9bqG1rnKI5/QOcK6tKJkjZxGe2Ew3BM
cCQkbimRjC4YPl/pK5HLmMKiR21+KN7za63uH8pGyzPsZpx2VmINq2aFXE1NqIUyS0/MTUqZ72JE
wuFNg7hpnbGz3x47m2BH+9r6VXUVB3hWjnDlxdkl/86yKk31jlGWVMzVyUoolhfcQC/fA6BhUBo+
x9PqJH1yeO83g5ZQpsutcRi5LgwWE0Ad3VeoEubUsoTaH0WsanLt8N4xkjbXLwaaPJgOeH+t00MG
OP+/szVcRISV1aUuURw/jcE3EZmmlYkbrpSFR0D5lLqBYPHd3d2a1jhJ5v8JjMxbpjEsSD+7aF4S
ugWmQlercJiwBYZ8QnQY7bJg/yN6hS6mXhoCxkieDnch9AsMOb8w2uCuq4ppAgiLcChVYRxsfIe7
G/+eKTkSBFig+SV7THllt3LmR0BDAkHTnZ5nSzA7pMqSt7uNKsZhjx7vs1xsTvnOVxd3alNbK58R
htmcqVpN8mjLGgPm8Lq/WSDBhAlPf/j1b3lfAkR7olR1uVeR+ntDx0z65PUg2d8NbheKd5jn+QkB
sqLFF1Nr/0ihnA0T6CmlrcX0+6RqUFhXzBeWLdIX5AUcQy1IocQrd86UMciJn6RUWNlbUWQAgSeJ
vz8ZsSkQyGko6d2pdytzBGYnICiDLkIr5EFlfHavGF7Q8CiSfnWUFWmALFmSNrDd62jdzjuOImS9
Z1naixRtVx9fnyYtdep0N4Pi5iClweslkQwihTBf0MkuMW/lgiPUAXgoDeMuBj015wlLX9bwfix+
jtL3NPLjfAmeSw9fSmgs1+d3MVnyUzaXOVr2oN/x+EmwgsUiXzxS1Zj+ukFC2a9xmzuhtzN+pu5V
OCQDnAr7UFZvWwpxl8mZmorZL+0QtCqGfeE9AsrkiinW4M2YLarTdr+msswo/R1SmdKBi6aoM07E
wsx+bJqiXAGFH9+SjkvNAV6S019Zia5Bpp7xstI7rt2QQd6Fhe6iFUXLI/dDFpSBDtupoKfZStJ1
mFT1fsj6GPrXAXGJ++jdPqtvNoWFqsQJj0ywJB0mx26bYISES1/CRSEykn4a6u9nCpLmzCo65ylS
H9x3S9qeVqPM9reWYxdQizMiVawt8joPBpq5QnDuLaQYIEXIC5u9Adgl/ShNGY+a2w/ZkKwN0gFv
kzFyNbLfVYe/LGaErd0ZYClGHy5NR5IfD6nkNWAwQSkBLbo69zoVBqOFeDz7G560TX9kmnp80LiQ
f2f1gi7He2S1N9ktgPkU3vm4Do9Avw4kFQ5wOmVL3ZkXuXNeJmol8AW0cL7mo2rOdpT+z1KXWvs3
Ao8W4/hadylhZfZkHHmrHf/979KfGJw6MyMuLMjCZDIME37gRt9MkgkQFeadd4VCZhIYvHJJjCTw
co67C5A//uFlhXGrBCaqTDFYzND0DfAjS5BXwgXFoyWDqvG9SQsSXkSF0oynOl/PYKhu8/GOK/7Y
/+oP5outvROPr+UbbSasYoQ7vC+68JYIiWQiYziGpEwzQas1iVLRUNkbKoQ51BzKhHReDnDprDFQ
fc/bFOyucTZag/6LGQ26Mne3oqGJrhaikJ+FbM9fDUOsz/JSOkNuRre16/KXF8kDz3SnI77F+Bo/
V7pxM3sySyok+CjdAYsLyKpMCNYLu0eOWbQr94ZKSxW3hD9DMd2bDvie2bftylBTEbNof7IxJn3J
dSzV/kQsL+je84g+I9L0dxDPqINRWTDkGWcKc4j5NWSvi63nfkdT5RbdSGbA5w0oUcD8YeX6zVTJ
e7liqEn/kYZUSDh3RLLAkGAmEVL7tYub3KWBi7LzrI1z8RIvHLC9xVFWqB896gBGnKtjBAeDjfWD
5/K938Uc8gDrbZufRw0uIiAuDSCuC0lcGUu3dFp5D/k30P2RE7zvEFz+Sa7TY9XyC6AHcIHjvPK+
6wkzA6ZbyldyZtmTUa7tPT8cqOAi+Phm4XWjOeJR8goV42CNnfzoSGrQTdJDNZOwHd+u8m/XPc5q
1Adth2Rs67eUclc2O6qgAFn0IVEbHzwACqFyU3RWesgtzR83hiK9BRV2pARW+tZMSlQ1FAEgl3Co
+0qwTqnTpAUF+2873x4nO7oGPv/YvqVPgj2PIA3pLGgrEHd2LT3PJuTcmfzGSd6g40eAGUG6T15G
eSFRF9+fg8NA0OgbIda1c+oUbcjaLuHb/r5sdPXRU1gi78JdlzXSLhzT9oHCZL543bevVOgUvOOt
WZSXSHTndsWshNTWULepnzfrxW2VbaPyJdhgsy0q9kuS8nKGLqPPsl/fa3+iw0hYVYgBSDSXzAYI
uDq/hYWXPZe0MyMi0DJ5lfwXoM9EeWjI+nNqeqlkJBhP4IJIXeZ7z20ur9K+4uu2s0AmY4lqswRC
zQh/0wPqfSLm2nN77sS/h1jvLl7XqOjl6b39XR70baH4ltsn4ilTkJ/s6npljKJaF5NN0cysTmxV
QeYlRyZTm3DheoP1dRi4HcS+MU7/tjWB53O8VFy+4NXl0AvkmlAukQrqhCnUyBsKRW2Uyf6xu8CV
dnVQuLFrEPxQ0grHfenBjbrGTD6u3dN5vyLIIxcSWtztYIehUe8sauAB7Pjo8WvHYgks/rYOhkEI
4VqHbs6AKXDxLkVcJj4T1gYRau9liymKbGBo/x2xqF1FNGTIx0pXpxQQ34yop9/zJYj6boCGnmJn
DC4NUYxtJPKh0odP7hBv2xqrW5JCHD68ahvUhSt7FKrJJq0LJVtO9RQDgK1gey2sfWvysHmb5sxS
AT+vXrpKDkDV50RKE+1TM8MKhrcG9+gvJSS9nchKAKa/r6jXhP/979J+fFBWFQiy/3z+3J+RcWaq
zaFaK6k89fFcbybwDuzggE5iy0D07BPV6D3iRzl+/+2Q1grH7QouiLM0B7U6IKTaD76iUYrbwjVn
WN7y5lHgcnl10s+NUNWCckK6ENPLZBU7YF28A0skuC4gRwqX4wO5l5DR6F2Jggh5csjl8aGmFh1I
+/kM5tkSZXsowrEBobEZKxCFa8pcVFlPmwaGu3/kZSKliU0dYEhp6Q7QTOh61UodBtb9cFyM3gfQ
mrxmww005IcRkH6s6iZ3JN0B6IBbMQhK93TNFOcciIe78gUwKKEUSkQLIcCANKsSRP/4Pbn9qvsT
kqZhcC7/JZe/+ZCM2DNUBnIKD7SiRv/e5FvQRXj3kxfa+xIklH5ykp4TXG/esK6XSGp3hj0PgnBg
bRXzjhMhDkqtoEYj+pufGik5M/HmGMDzhfYe5NP6aMIr3rkYzDjD3DxZrRxb6aXd32AvAf0bVIv9
9MUf7nEJ97t8a34klTRpFqOVYlnOxs9avkWd39mNuCFPl7ya+07jyiC3gkd3pSSQgICZfF4hv5tI
2D8pvS8YSP2M7mRFTVo2j3KYIWTiUR7TGqhpkBgJOkzpaOq4WWVIvoVVxxQpixGqUglx1oVNhBcU
aLki5Z5w2PRVvO+qO7n4RMNGt878vyOeY0+PTsiHUV+PjmakocdJU0NGPKZ0pIi4D+HUWyn8iFiP
AUJ/3ucPxiT3D//ZlNwPShcRHXGC1JOghBJeD5V0WBomArBZhtcWDyNihIw84vd13rC41OTvekkr
Y0FPTH/aSG3EdWK/V1FND4HDtiWnClZHHVUa0zU3/4wKnm9H7vcCa2eEL1VPVhiYcq8uLtpyBchH
Tu4mfMdsohSjzBa/vOi2sb+ejriTMrCvMbXl23ufBUHTaqPX8ku8S9U3GYP+mdInYybJi+T7RnXG
hJrwhS0joLUo88RLzwyGDfLjsurmpgEG0/mRdivSoj1i/to/x9sl27yJ9SFAtRjCEH2tufOgeBA0
pDdKydPJWFg9q6cF3TzklcdkcT+tpOSeBMugyXG79r0TK7b9aawOjkrzt8UgCe0/k4k/zQac/rl2
eqze5yOtV/AynhS9qEVs4YHyu8MyOKSvr0OOgQNWF4zDAnA6IOV8+yRgfEPYG1UG3HighpXzzQuE
XvNoAnvgR8ZXsfGIt4EWqwELgWIKGeolSUG/mObJ3Fy8N/+iAw3gBnG9fn3yI+n8YAB2PQfGx+tJ
QmqU+GLugi65OS6/sAbABGcUl/g1n05HyFkjktBmfWB+tvS+0pFIdDllkIV4tsMKX7KlXGVgCepB
JZXPeJyEzXW5DMiM20h+p0H44xM5XJv6QdH8rrHkxBkt+vogVWz+MrmYWva4gaT5jxm/GN4X1zgs
kboVx7IipnL7saZBdKPUtTu8o1TQkY1rWAzvc0BJcI/TM9o/ZoSmwvUl1b7l54R1xBipsOFznWVk
PTpbncyUTr8OjDj1UPVfZYnN8vJxofXfFYGAsPeZ4VxSkWyYBEyVlXWn1cVAD8G4o9X1UGFwyLEV
B8QHR6o5mP2H8wSrK7IfSAuhRZy22LOu6ilpd+XtdFMvHi3FnbC3o+H89sRpVgVKdCbdkKYfp25E
exILp3rL/WB2fZfqyrDlBH/CvbrEXXBwXliujsz6WYI1Z0ad9pUUZCCwFN+iWVdx5QBNzpLI4fiv
3+m08XTMMnupKabPRWAuxDOiTrz2sCcAWqvigbmuH73Wz7I27lr/KdGtaOP/J257Zai0hhVsi8/c
+bDM4fg8Oj0vgO2UoNdbi9clSx47W6oQmuxsZ1sKnyqLHEsXPeUmtO1a1PPtTa9qOsBQ1UBB8dZX
aUDJr+sLozYJWDS7+vlGzrIARgPvdVGN00iY74jXvJPxQikS0feocrYg+lczABoshEnURDmkLoKm
SV0zVF1YfxPppCQf4eqarhsNMD6uUXADX0pM6Kf2/raWUvjD3V939N8Gm+M+IMVTZT/e+V9/q6sx
wVw9XVawm2PqOuK37tvjnf/5ySRruQiKI9AxDO/lSZAp+Lz7Le3wTT2n9jRdqOpFkC8MbqD7w4gv
VzGv2y/kY/egfmSEs5TviTRjSpLNRRbXfPSznvoTxUjP8IlpudvCrsWh2Me1dZxEXkVmmhwtJmKJ
a0gnKKFEr+c0Ey5+mAV0lykh9zBU6znZ7UNDZHzEf0DGa5k0UYj7Q0dbMZpCjszrVFeM0tA3p4/t
w+RSueTV3do2UTs2c9qICOe8ODWkgHLOJewy2DIiZgp1HvsIC/y7vcoWEsrpacjfff0vx/mY9Wbi
0rlw7V9FZ0baBvq+tcRPxmIqtpv/1ed7jsRX19K2+YC0+epayya8rkHCA/jN8sP479juDjDr0hcY
g0BUSI8E1RaCsG4B39QLb/a9f+VvdTNcmGERi63vwpRdZX8OVD37S0f455kAw5UDQYtZf46Q4Gg8
04t1JHPVesnvlTYo91tfYoFBbwxcRWrdwc2q/T0DZNWLjhMjqKsFxvd6md8doCSTglExiVCCapsE
yz11vKT2MFsG7Vb8pYzN/9wjXeqwEGjJxpcV3C1fQ0U4uV5M6P79q2zW4vgs8v6MYDigROBnBOCq
v88mqFJtqCdhJOTBmum+DGyitBg4zONBKPC4SPX/dWMgkCZIcA2IJwj3EFF/ehMKqwyvmsMEj+BJ
UWAIy0Q77piBmn5dg2TQtkb9Wl+7EuWFoINQEHedhNXPg0X1GxkTpZWiF7x7JcbQmj25CCyGq8cA
ox7M3mvFhhV10c5/PAogWyNXVm9i7DHcScklNUTqYkEfCwSGfndLIHUywJwsH0Rc9F0V9LVA1FZf
+yKa4Nk7rQJ5X/oBIwueFakKealMRWj/A7WUMn3Kzx1Zv1lgRuqiCIYO85W15hRTkQ0yXGMGjFva
lHbFRBmsdm88Waz57ihYXdwpPYZ36N1c3bL3BddK7ZGqoe+CpSM6YQ91Gd0sPFkYc4MZrx4wj5Od
EYip2e3EEKjQpa2oTYhDDYnYBxpttQrgCV+wD+FimmStqdR5cCtnEAjF3vBBdwj4mlK0964nbBC3
FwGUp86cRJwsI0698PlfkullTrKKClScxQCaztjniM9I9g1xVEyHgCF4BtPbI7FeWND8IHuXoXJr
uu160W+pr2QjzuaknWjUhmA3EV1qS4hIYjrfWvCwQkf/oX7lXcks51Eyfqze1n79bU2xTdUgYU83
QC4eX/f09DbKTx7qBe9Oh8zIeQce188fXxggSio+UV8xQpG0u4gvrnejaI2kKC7zzcr4sl65omfY
fUC43xfNKckz3gAkpxJ7j3ewlv1cpG3GFt9aSg+O3oH+XN1U6O20BIKDTkCaafageQu5TuEzOU9o
jrwzykusIELf7njYWSKLyjCqgsKWUnFmIsMh4IeJQs0fDInYCJW5LgkNV1hqIouvQRrZC9aTY7rN
tprl/sZ/eMBCJXiu3A+bMr7shUbziCcnD5xvDqiYko5iEW+MuGuuK0cjnwF/XejvhCwzS1BiP4h8
r5rQ1e/bHy5oS3OlMBJ+fhz8TKbcih5idXJigKkAbf8Y9bkHKq7J7XhmEzHPtYo0Z47tL0gW396F
IXmSJTSdUjzs3Cjr0pQEffg0qIunHibiMr/W/TbrtOLEgLElKA6lhBHhB/va3IaVvKXKWS/tnitN
uEyTU5IEfZRMnB3iequoywmXNEnOrCb6+Dmsnnccqs1ZLzzNFO0NiMbi1gMvOqH/VpvilN7WKxpI
VNG/T5PxNrZQh1VGmxIjQCwSPvSBtKZyNrxVs5nH2yCqIdQtQTGgxcZAK8ILS+q7EJ5QZLAqPWl+
x/6W3RIB33eK+Q4gZGTWUpw2z3+F24/3PEbf7UQ/T+g36LKelqRa69Obu52S76cdOGR43kM7Dyb/
G9SLqvbMCKPxrOA7EUMvG8uVqhfO4blQ7ZnPoAriZobR9pD2CCzYl4p+mYRCG7sbL/smyYyn4cW0
a/RwjlR31JbFG8BzqahbDHnXslnV1l2kYiUyyDdyoTBFAySUpoNBTnQXDTEemk0BrZLlcFrQevUx
/u5sNzihstPnLWjl/I9Y9YEPYu1LntKfxYOBNkuFVNG1Aao3aGWNegrpuwxvjgHEuawIo/tPf8yE
GrmO9CzDU2S7SWF7KO5CMZHWvvGGQHuFxGTpzYDKg9CknOtW1y2XelvjPY+0rYRAbPNO7Lc871Ca
L9q+iDmewpPyQ1YZmqgnODz2r3ogc59YZsCEB7QKMjgonvPfrl4ZaK8r64tB+n0aNMs2kGHKl8A+
i4vXQtkplpc1zIPc1cVM+2NranIDy+m61OfVSIooPgFXDBsl3pLoSh7YJ7jas3YFFOrAq9V6u+Sg
TF1vKRAStcVMWU/cX2Qw+BhXmXL+Ua2qhArtmqAbcLAQkltJN1XNeZr06Ys0L5rJ12Ag5I2ZrDAO
iwLBzZpTl6AHQNAqtQyFszDvnT/5U8K0/fGwWRPKvdUu6tW9aI79D7eqnWRc1x+7aX9wRDaJgbLI
LlfnLub1jLEGe+aJxof2udkMFZfgVqMzLcspaSbsKeio36HEg19fAAwXxiucoZqbXQTGfSBpI6mS
HyuldP99fsI6xErjTzlzDoU3nR7vuwzZCYcN/hAkmsWf21kqpFm6J5iDkd8qMVcf62N6NKo5+F0+
WsS7G8GNuIQFIh3AiBiYTJphUlPiImfhvzRUcOyNQ/rUq1j1kebwCidoSUSmEIOnbVA380FbUSOr
/FvqwlO9JfxodqgvJdmHLGpjdUY8QVpfeDW+OsnT+veHMGL+oub+fUvabJU9irgoZ/6pej2yD0Bv
8sRApmnSOBALt1nFKDPxnQ74szyqxQxxXPbsJ/gOPytsZnm+GAGlBG5382rMFOyngLu4+dzNSsa6
/7c4lSwIw5Ud0dX9CH9GXNN1/KTdoXa+SBTACih3/vuf8CL+aowmX78vUewRVeWZOLR4DaA1sNIt
BleaXenEBVEsf/s22157HFwiHeipYl8Y4gUseoXLfvv2MEzTErnpkQBoLPp2EgSNPlhI4rT9oa+T
85B5X+aA0fzsXwvENsITzng5wqrOBNVhoHuKSmU/9vFnYpyCa4zhKU/mP6uJDYyStFRBLwL/SKaB
+oc+4Tn/kK68qkPM2QR0ZcGZb2qbxPjIVfgOpl+av1nXjfkhYtWJFz4PdUokAQAY3Z6b2ewEBQX6
uN5Ie74BLc16FGcB+BbwebFsMUZ4yApoACVm14dMjjxrFtTIMsBsGsINZRyOm4GrCl9uMN/wdGOA
wK5zJcGTEszY7j2VWQRn9rM0xK3zxQXKViBfZXl5ecS6BWQrCenZOURv5vx5jLzkIHw7n3S+Avs7
UKbagm3YUmldLSYKRdKDyaMU5i6ev6Ebl+vnO5aZy0Arf7SaEmyjJOPu9tZzcxjkCDG/tX+7Lgya
nYR5mrXf2cuaiB6gBytV8zyMecaN1kfV7sFH0R0qA1q0GzeotaKjgqJuobvxBe516oyOfRUwaULS
yoKAz5G0ncDnrL7ZoU0uk0XugI0e3/rrW+ojAD8nMQXNqmV1kMOKRGEIfFQXp/OSqI6MfTpkDkRy
zrbhmetEhBFMwjBfl3UkFicplR312CIlxGGVz3lMPSpV//KhweJ3WIuQJ/uUhDUUg7spv87Qijg8
QUYqmdAq/jqb/Gev/RaEZQVxD6rshs+RK7RZ3m6EbwMUJcgVKgerce1SXxm+ULSmgF6Ly9ih+mbE
PpGYcIIEzTzK3SjlJPcpGXjRIGGpYaGPPmOE4cW1aEl+yA7SJ74O0ui3yb6VxljnXGeNEdHpSyyB
2baXPG9sd9jPX88wd/tt4OSkqus7PH+6eTi4rWJ5ko8bxtEZMMbhCu0d5o4QL+JY7C06662UK2DS
kHXu84PGhcO2WhVjz03t5o6h45nwjOGmabR8mwBy+oE4P1iEo7u7zaN6CZMB2Wrr7dv4zy2Kza1k
dPs1J3IJCO4DFGrHBK7Bjh1UNaD8pn6+Ve7qfdF2spqtcTFK2I4KuSMN/+csYu8db13XRUbtb1uM
OEbCmkr8Wv1/onPOd0j+j/5dV/8FUesj6othw65x5nGO24okVAoSCvaB1LjEJCQRAxhO3FqVouRv
Hvbsvqvohb3PLOsandSixS8N3X5/A8jT+3IzBlyRjezbYwQRYqR0j+1asvhU3mJrad+SB0HwQvVa
WAW8KdKGmKWCUFCFZwZzYQ7dzFmrC5okmatqdI51UImAWneTeP75mqUUjHoyXZch9AzW5jTqUBVP
ApvTBLycQhzYkhgMywAEZsoPVzy5uIoxZMv1poSX983Cxa6dClewFUkaoB8nsqFp5jw33x4JLpof
DpCZtkyiQ6dahOM2MFOUuJgboC+R78lzmIUsRiMq8Gkwq3T37u70OVBBU7uAWcE/rBtlfLAJTq+W
EBwX/o3/79Rh3PtHT5GRHchvYwHel2VKfeaRZaTPelyJP4qOQNBDbS5rY1+Hb0ScH6kgkRMUNC1l
ST88saPwCD5A83WdBxdX6OQ/c6d78fhzWon+y6FDWTuZgC+kwXVEZv4OrA2QOvLaP88cbmv9/1Yn
JXdhRTXjLogHSNEhzg2klfFHO9yvz24NWG3hX+O6f8O0Wj1yZrHomLeoKwswpWBvRmEKwg3sGnt8
Amsgjn03edtE9JyXzgnisE0ipp97Wm1EPvWtqHIlVTfnT2znzGo8rpOEeMOPn7cLz1Gn4XUnfwVZ
1gmecC3Fl8lVxUj5yYCravtnPvCiEsGdRXz3f8jbsdi2Qv3GAImKEg6w4Xg6Q4SxmhTawJrMW+RJ
QC0RHl+owMYIDP80PzKfNhAFyjySbYr4/mhBng5gEa7/BKfcitwuQ3TGDzdEOPNbB2DN4Av9jtwD
2n9qzx+7Oi99MOoXP2b6GkXpPGTOj10bgkk9/0xmKkrs/BhsRe+XFKdW9+2RkGBz7kwsqlUlvl30
2gH+Md05yOhqXWYJTNdgq4upUDqrjlqexqXopWzJnJY8vLfA2g38W3+CEp5zc9I5coSyD2nay62m
SXkSb63wVKFGRsgqN4uj5hgWH7CWbCz5x98gUVUcCLGg6WY7TV+/HTPsLpitPxqKR2xIC6zdi86T
G2u89VMeTD1e70C2SaEnujR1GRaDxfpjW6ltJg8BFqSreTWDDIKP4fXVGuAHaUwdNkQy9wi+xHSW
U0b4ujrADgtW6C5S/I9oCp/aiL4wXFEAPTBXgjEFpNsBYejb0F9SLzCbjj3dfTLoJIkckhwBSpmc
9cuq+Rp61BszBrzLZyTC7i17AZz1JXzq/b0QkwX35qMQQqSwaeFeuGM0bhMOp5ojwDfugdDS3b9v
i0DzatSLNpWLJlJHyW82O3lkD6BWwKNMacKzNob5RqbNWts0xa5t4LT4WtDkUDnO5vIcPCwcifk0
LSMujmNvXFFTjFxVzOQUzTeoGsJFCgiL6E0nXfE+D4ydB/WFMQ+Wk/F0tVxXQxPujna1QzsZuzy9
i3lxsdK4vxVWAui9wICt3uQf7jmWfGEcrCMGlbsQ/a75TNyWqdzsHYD2IEhNiXA130IZ59ZaA85v
kC9/zuwCM9TfpIjxVIaOQ+n/U4Vp6VNQuibazopc44mJSg9xhBxXu4tnk5rokOfAKSEQalKJaC4R
TMRywaEYE2lJFawDaZacmU1A5Ulx+KBMAav9MmN8fe56Bod57erYUCEhv1SWODWaBFGAibPD3jBs
W6JgJONE/rEkIxxkshyxqemchc0aoHnDTM4PQLpePYJ3koDNmu24nhYYsqiXwyvJyrtKfOV4r+z/
sH05BKd9GbmC0D18yxxmBQrOpFtBKweZKWbPFunS/K6bpPMSXHsJWXTHwtL1aOeRsaN/sx4P+3RL
CC/OOuEnwNP9dOMg094DM0HUN39kcY5U6dNxCliQmdVgxYgk9QkBkb6HfVWaSQJgex2wIVeJLr1N
YsKjCDM1RPc2gdomYOdb/9+rXu/zqcLeu+aRFTpEjYsST5xrYzJWMh43X1CLz/R0ARcvnECellvC
stKjv4iGSNVadI4sfRorhLf5qmHZP4Oa+damAuyogAU1+yWYREeHeIaADuflqGkN/aoEzpk3b5wf
I+tmhn97MULZUTKCMP1w2YudPaXr3o0+7EnB8dhJeAMDiRVMYWoFF6JM1oVvRKJAP6/zPcof4Mnr
jrQSNg0nfTQwrKMhJdbcmhjigzr1dgslxjYBjOy1rOZgFWCzjhgk4uov0bgynO7vz5672fED/nQ4
SF5QUP9s8otwO6bJuzUmJ25/rDqonei5RUPyjiEFV26kwZGpgVA3Vr4aHFAULf7zd0K77gULugnu
aYl7NKBji8ov2MawGiy/Kkc+rwjbDHT9fpZMITwDj8uOAqYiac/W5k9/WGdj45wKU83Zy2KsPxl4
HPjLKOhrObYzEkAC2GfV7meNikOuH1bOqvGMuE/zLK/AW/492ey9KyD23SqNC7Q5WdJaS+6ILwCr
48age3pU+SaJAeJ6vB0ZetdRR+8zzft2+NbQQLF4aDH3sdAgaL6OswuzVJM9+Lsjk7mN24p/2Ub/
ovrtwwIEVs48EA8Q7nhVzDi6deLKoacVwsw9/RAyq4hvhAolqmY/N5jZDCinhwqUjYE9rsyKmojR
/x0xeYi0inlwSZLuRAXD0/2wk2aYCUYuDqxl9a+FlK0tANlEcCSapsBJt0yKfI9Xm0Qb3RX2AE0P
Oom+yfwJHIOoo/YFdEu1g6rk+6JIgV4bxKjjCLOHXeEAfA0ZfC++4qCjyKKbX2zig0W0QOfL5wBb
ZGIRzFuh6ik3mgZEPbJERGdWGm9fOMnaqHEMun0E7n/SgkZm1zlec0cdWUPtAuyGEi9uIDVi98ZZ
YgMY+jbSa2ldyZ5LI0I4mADRHYFJMgaDVj3JSTM7QS/wWOQqSTFblFwGgMxDaTVQAeHKkPisYUC8
JRtkfeklo7uQ8QcHYse5YQTBZ+UPnMbg/23vUiTRY2MlY7O6lWL6pAe36wWRZjcaiS8vz17X0x8S
x5dkYp43f8IHVeCq4t3QQ3kSqwbVnCnO6fKTKxTLCoGmXRFPXhVGDqJx5NG1+FxyOlb6QTdL0EiA
/4JLiH5X0vTUxJirUGWd28/M6PkEqlW3S1Ri3iOX0A67IT3fOttvzlJnRkcgfFskImAH61I6BRzJ
1QGPOQfLjiE/MoZbV8t3SF32zIQeI8grRVzOuUwogi6RIvz7KyMqV+wA0PC3nw2aVeShPEvWxbEb
/LkZt41inGvKBVFL6F7ikxCWq4ql7YMnT+rfYpVpbKfsQzlUHc6+cfUSS6A0LYk=
`protect end_protected
