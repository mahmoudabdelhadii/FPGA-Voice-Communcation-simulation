��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���/�����Cc��<Nb��.�x{�>��0����=�����=8RLG�h+OLزV����ݗ�@��&�K��4cbXu�6@A��?��I�=��O�s=���
�S�i\��D���d3�q	��9/�I�w`W?ދ�S"K7��5�,l��C���
@E=D��!
����荾Z�V�h��c,Dt��&�����]4w9K_9O�=l�uE�w����[R�\�zÚ�-J�$����åCj�[�
����T=���K���h�����,������#�z~��?�G���B�~֨1)��k��yq�$/ju�YA9��SX�{@��mWt������w�F��r���������O)�mC�&�����$��^_��|�����=������A���_"�s���50��-�ݡ��kVE~�cu��'Ah%�����v2ݲK:|�g���7/��=Q�u�~��qC���
qSa�a�n�m(�]�h-�FK�]�Z<��K�b�s��'�����C$Yכֿ��h|�[@lXJ�*Qm?�аR��(�v�vlr�j)ڦ��0p�s�bv��jy�-����(��N�vהS��Y�n)!��\|9��;#�o:�#��9|TWL��L2=�'���$ƫ���19�?�:H�A���T秧���,rJ$�p}�a�ڡ�rn#9���~�1e�[e���!������{�T�7���O�z�������쉎�<o�j��D�7��lS�ƃ���F�V�:¦?�,�:4I~P�o6����2
�ԫ�#��G롔�qH���'> x������>I�nN1.�yφ�V�ǹW�)��	�3���k��c�Rw�buRA�8����\��L+p����rw3v�FF��8��Y��8p��s3jL&���9>��y�(r�I)ռ�I�|���Ք�������be�;��5���4����;�4�W��K;'�-G�#�����*����uA~���Cмojٳw�A�ڣ�M��3�n��E�BW�����V���4tDt�5<��=m�h�gX|
E�t�Y��~�Q�j������:�I�����韰p������ikp�/�4��Y9���i DW�#��cl3U�Ty��PH��3���a;�%�ë�!nd�(X0T���`B��2&\��D�c��Q2���i-����̄�Q'Db��Yg��g����E|s�+�J���	�8� ��`v�mH�H�vk�u\36�6�`r�L����̠%s"��|e��Rg'k]g����Z�Y�P��:�qEr���P�S�p��+k6(&�bU�Y*�as�sr��H/�_������y������]7�OB69}L�(�cc��Uٷ�QH!��S��~a�:��+�e(�l��,��*߹�t<Pw8�i�'�d���H��5�7�we�!����2SxG���V(��(��{��n��.O/���[lb�l/�n{#aG�vr+����Uv�,�?xq�����|@���p@2-�j �'��U���3��
�?7=�����o�rl��!GMkK`�Ů��O;�Ӑ�p���I4H(�	.���ӯ���%2Τ���O�I�T�ۥZ�"�lD�;�,���ۓ��~^��s�����$�^����Q��d�zRӫ7K��xl��um$�զ���|���_�3��R�����FQF'���m(���H. j��8����$gA����q8:�+�$(B����%m�e���w�0���0'��e�3����r$�jP3z�P���.�=�P�խ��:6�P���/� J�H�9�e�U|���=;W�'ܵO=L_|8c��L��nO��lK$��փ�F˰�s��,�g��xw'1.���C��>����>�u�w��8�xc��"� �\ArVƭ�z�~TfH�˔�1y�ڷ_|/�������F)@ynܫkl=Y��E�]!{avW&<תSѡ�1�<�:��N
c4�Ҿ��g�r��?��[pTR�5����[����^��,?��wV?1���v��'�Kj; K  �GP`{k�D�����T*E-u@@F�"xF��{���#� �H�݊��+��D�|9��0�6ޅ���F[T,H����YƁ���ۇ��]���?.�9S���Z;������m�i�%eG�x�,��+���mZV�����/��:��̛�A�W�O�স���>x��k��7+-�|V��\OV��]�ⳬ��gG��~�e�3G�p(V�qwz>����zm{�I'G>�I�LY1�ѳ,M�#�I�%�cZ���Q��E������k�.\�W�D��(������
x�Oz� ��2)*<B���ͧ>*�@h��a�0��Rff�[3*g5�ֆm�3p�[;�܌�u����KB^�7����r�s�����挏BE�;�a��\�)�_^���8_���&���e>*����[*���6u\_,'xW�	���T��/�}���Ȕ�^�f��>�E��'ٶ��{�ν��B��y�7^ś�h�Jʻ-򗙌f�������ڴ������V�h�����p�s�WD&�O���:�n��̽�������t�Ī �GƮ��;�2��N�Ѩ���/Ju����ػiw����<Fa��c�_U�
D�����5&�5)��[�l��Z9/Pm����8�6	!;a^\.1�	n�9�g�
p�M<Z+���^1~
#Y���O.���R9(�����:n!q:�nsF*�Bɤ���P�֏����@�!j
����*��=s�9�`Vt S��	*Ӈ��w`�3��%n�����C�J.��^A���~�Z����:���%��l���w��\�z�]�n���#�Du5p����j�Z]����+YaG7���a{n�M?��t��+s����j���姷���E%B�� 3ui�z~SBS��2l���[�E)��:ļ@���3"�������},�z�a70+�	��W�Jg�i,=�L9�
l�U� �ݾ.SE��x8ϼ{�#��s����=2Lcu�mՂW�Q6����ͅw�5�UW����V	G"bU�<���$9C� H�;�hi�(x����qlt��(����5�4`^9��.�}�H1� s�X�)2l�	�n��A��\��4��K.�PMp���r�r�)�w�o��:�/��01`�Y�ʸ<������(a`���L%�nՎ�C��	���,��z�u���)� o�C/A7X H���6�1Ї,���)���䄳�y����`m����|�Ke�(�v�,�[�ᰙ���4�:�=�~��4й��P/�X��ׄ��O�.8�8+|j�������҉P%κ��z�C���V����4���BO���J��~s3��3w���xj�b��
!��g�j�v�$C,`�y�ѿ