��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���/�����Cc��<Nb��.�x{�>��0����=�����=8RLG�h+OLزV����ݗ�@��&�K��4cbXu�6@A��?��I�=��O�s=���
�S�i\��D���d3�q	��9/�I�w`W?ދ�S"K7��5�,l��C���
@E=D��!
����荾Z�V�h��c,Dt��&�����]4w9K_9O�=l�uE�w����[R�\�zÚ�-J�$����åCj�[�
����T=���K���h�����,������#�z~��?�G���B�~֨1)��k��yq�$/ju�YA9��SX�{@��mWt������w�F��r���������O)�mC�&�����$��^_��|�����=������A���_"�s���50��-�ݡ��kVE~�cu��'Ah%�����v2ݲK:|�g���7/��=Q�u�~��qC���
qSa�a�n�m(�]�h-�FK�]�Z<��K�b�s��'�����C$Yכֿ��h|�[@lXJ�*Qm?�аR��(�v�vlr�j)ڦ��0p�s�bv��jy�-����(��N�vהS��Y�n)!��\|9��;#�o:�#��9|TWL��L2=�'���$ƫ���19�?�:H�A���T秧���,rJ$�p}�a�ڡ�rn#9���~�1e�[e���!������{�T�7���O�z�������쉎�<o�j��D�7��lS�ƃ���F�V�:¦?�,�:4I~P�o6����2
�ԫ�#��G롔�qH���'> x������>I�nN1.�yφ�V�ǹW�)��	�3���k��c�Rw�buRA�8����\��L+p����rw3v�FF��8��Y��8p��s3jL&���9>��y�(r�I)ռ�����LEe/��5mJ��V�����C�Һ���� ��}�q�����쪦qe��й|i�<�iC��U�1>��<	D��;ns���"�;��ݓ�wD[�Ŭ�?�f-ߠ�m(aѓ��T� ���c�&��ڰ엡�o�a��e���&�>�lfd��&�F��LkP�!����g��潲(g���ބ)_�k�"�}ɯX}�^*�Fx��7=[��jƢ��q��;[����řZFP�z�_e\I�|P��؂�v��Q� ��&6��CwoQt1�VX��*��-6F��Az����I�$�+zn��(g��I2��8��A�/����k�=��=�M�/;8p��߬�t� R{�3��Ӛ��o�{����NbE4��&�Y��IE]dqw����3�������8)5���b�x���R�v�R��oc�f(�t,��TF���6���c*�#� 0�T[Y�]�1�W0�����(�'��xѭW
�����_�	��Px��H��F�Z]�]�5����+���Y,���[/d�\���̽�W��q�������'\M��u���� 4�&����vfd�}{������*<E"���#u��)�R(�8F)"��B�/!3V��m�.w�y���	<�q��-X�y6��Jr60�2�ʇ��(4�) ��Ծ���k	-�����Y����?-ɺ-���#:1s�PR;V}�DM��o�W�~-:
\�0&t3c��cm�YeX�˄A�o�Ǌ090YΨ��� `'w�q�M��Wۯc�h��\����aߘE�1�w�Q�]��9����.Ԥ|Od�1]I�PP��awH�4F�(%ǚ���W��}��.�NI?a�ƣ~$%% ���������q��z����	�����G����a}�2�ˤ�W�&�f��/���AV�(�9�{��1����@�^k�q�wW�nz�Of<ƞ�N�,�)N�h�ps��p"Sb^
��G�c3�%V��,����I&~�p+�- ���5�]A�6�*��+)��m��+6��$]�X�ñywT#��}6a�T^s2�Yz�����f!�A�5�c���[��LxT`��LɌP4A}��E3�YS�O�]�p����D�b��{!��럂�T��!����_ �yF�����/v�%QnA�JT!��� �.����t`��@YX>�"_�kR�G�ћ�M�CK�yb;�癪2.��C`yD��k1;�����/q�
38,�5����Q*�A�In�6�.�+X�HN"��t�.��xk�z�Ô/_`�.�呪�(!v��\��$��wm[�U�ξ*T�����w�+�*��c]�����c�v��T0a�A�Ԇ<��t���R�Z:vd��8�8�m�N�i[!n� ㈹���M�]�Zfc�.����lꔁ��6�w�.���-v/\�E �2�y�cK������L���������;�Xq���]��/˂*�G.�-ޅ�P.S��a�#��o�obe[MS�˻'�������tо������V�Q�������|QM����B�9�s)*���g�˟�����܎TCs�@+g��}>�F��Qᮔ����\�`]<V�-+)u�c��fi���d���X��uG�g����n�CJ#AD8ѽ�Y��Y9e�dK,	�-*O�CY)ܭ�{UI.�_��^�	��6�����:m�b���e�х@�+D�ٷG�9%!��67��!�d�R/="ɰ�>\J��9���;�"Sd���~9��x\n����+ȸR@/L��s��0w�S���'�7Nm����T�C�AF�@׿k���}��D�zt��ꭦ8�P����������*��2�Ӭ�Z�8�W�P8��iwr�v�L NY?� m�`)�s��Ŕ�B1�����1��i�f��1Aь"Z��t12KɆcǌ5¥t5λ=@�!�v�\p�m��E�`i0	-(���[��<�V�ن������N_�Hjv�jcO�Q�������<��)KU�O���ߖ�����4)�g86c4�'�Z\���6WΧ��d����V�\��Q_�����-���0��XS��x~Ob0%!pѺ�����.�:��d�����C�ϸ���[ũ��V�y,L�ϯ?�$���s:�a��)ɻ�Jp�4a
�|��>z��zl�P����/�c��������m�q����)�YI^��O�lp�꽨���+�Ab��Nsځ�u���ՊS�x2{1�*�h�Þ��ꊅM������.Cm�m�S�?������!����v� ���,����: J ��FWz�uP 54�B��W	��/�n3�y��r�
�$�g~���4���
& eC�7Sܧ�'�4s-.�:�(MO�� ��$��$�y�8 �豨��4}ϼɇ~�4=�@lf��wu�AzT� �ɗ^rۗ�$`i{t�l��N����G�-�z
&3�**�j��9no��F.q��<|]��e��7�9���
ǭ��&F��[�� �\�?Eo޶���U�s�B�҈�Qޕ<3bV�*�L��C_��� dF�"ȏ�'؄{�4�y��&�%����J3��.�h��2�S�l��o(���s��؃2���k�x����)jq�!j�0��r%Y��ݍu�WQ���Ė�0� ��Q&	<i��o6n�K����G]�R����"BzX�qIy���?X��Q�̅�&���c.�Ƹ��+�@pt���:Y#���L�uo�,q�<�ӵ`�쩗����>�!6�����M`�w"`p����hHyF�sO����G7�pȓ`o4�HØ��13?x::��Y��"�#`k��)�)N]�+�2/��ѝ����+���!k˞��4�A��:as�I*�I���[�Oq����Ng/�g��k���������!s�k�����j[S����9�y>���T�{|�S���i8&��� N:�2�.��8�%�m
=ً�Cr�\��Ol!�_si��sb3���!���.v��h�Y�����I�4L(x,�,��$�G��V+�
'�Q!?g0=[��5����r\j�s��� c���8�'\ o�2����4Z~�ِ�9�2���~��X����U�{N3PY�i�b�[1]UǦ����ER�d;���w���+�s1��S��~����(:�1�e�-���M����D�V Ղ��m�.��;�@�7V[:D
�e �������� Z�9����ꁽ��r�7�9�2I��2ANܶ=8~��hߞ���X5�"���eM�˱LqY��e$���
yqcP/�r�|�����q�9����H^΂Lx��2V>�SL\���#;�,�}ޜKli|yb����mcB�ć�	����(F��V]�s<X_%f_L~�C��L�BK��"&�(��S]�c��S,�چ�dx����8�;��D�28 /�t��Ҫ 9t�A��k����[�Dj��	�s-L}9^� @��۫ǣD�rW����'��>�Tǿ��	�t�=
��	Vg��z�qMg<�5��H�(�>���NO��
5y[��b��g�J��
�M��u�w��S?階�x�&����-n�O�t�\[MC'}�8#�_�_�4:G�k��-�ț���`�~-��,���p����c��r��D���{�BA1�߭�QRF���#= 2!X���̩w|��U}��2���3{�j�B�z��E��;&.p���Ez7���=A��'y�b-�7��%g:�W��cO��$<7VE�,AH���3�P�7��c�e�{�v�~����_U�iތ��hK��x����ܳ�SA¼�^��mc�	�ц�7mG@(
Dj�%̡;IT���ߋ�UZ@��dD��a��{������a(�TR=�m�[I��ҲVe�E���E��T�:Ԫ���6t߲����3�V����v��ǁ�)�{�V����t����א_������a����-"�Tls"��,|GT�6j��5?ϼ������C)����&�'�1��-}wĸ�`o��
�S��U/hG�t�����wJ>��r���h�л$9#�(ܟ�%Y+�V���2��g@�2�1$B� +2�T��Q))�̴x�.�!>���hhYQ*�{� Ն�q�z�I���-�-x2�h���{8����p��ڣh`�S�ئ���F(�~\z�Dk<)�la�ڜ�k-BڌԷڈ�)�Rܝ%�:~E�� ���7N�D%�.҉P��%�"��ߨ<��b^�4��n��L���(R'�M�
��ɻb�%ˠ�j�=%����h�*'�;cp!��v�CcϠ�'q�#�/`��U �?��vBm����c�)-�MK�1D���*G��2`����4�}�9r2��2�U���)TB�wh�T<ȋ'9F�EL����-�n%��Cm*/i,-(�4�r/L��yr;[��N��vF
%���u,ޓY��lIj�Tຼ�G���H x��e�qW�bdq��T�Q)J�sb�0w\��\KW0�M�M�}J%�]�A�ʥk^�  Q�E	�HKFR��T�`ʠ�r�jw�cf+n�5��ց7:�8k�6-?�yAQa�h��sr��\m-B�c�pw����Օ�E���̩���ؠ�jaHbn��Գ%�)v��k���y�;.���'H��e,������Zu��:`C�8�t�@��{Q{��b���J:�����+͡��2��0!����.�&�Z�uG�����h���x�<7�O�Z񾭛	�N�=c[|����`R������mba��5���b�$(-�+���l�9�T�|�
(�!�c�����`_�AS@�Tz�h�	��I��}�`\�ә������I�cc��("G5'��)o���1����ڬMH�}�L������%I����:�ge���	��v����j5ad^e�<�9��n�\i-����'��R7��k�.A!�A�}�]}f�� ;�{���!
��Ǖ�	[@�ي1�䍕�0D���A��ѱ�e�O����i%�l�M])���ή#`q�9�[=���mᅧ����M\������|�4�P�����X|"��_�ΦI��Q��ͻ[��HrgIB	9骠�9���2C����v@��ʩd�C�{����K����������.�w0�3�L~08Ȏ̼f�����.
�[$h/$tWhz�~迈r���g~P�����]�ɉ����4>d֯S���`��Vb'0��[��6ho�e�V"��D�
@�6���������X��	�ض'M��ۉ�ah��R�&u�m�Ro�����U�����7�(h��;Y�j�Y��3pJ��l~���NȀ
BiX�$���Y*`{����v��t���}y����p�c�v��*9�f���a�TZ-l��#ED$֡'[�Q���\9��:g��sO�:��uV��uE4�k&u��r7�-|�dה�6x���-��f��+���i?Be/����Z��x��z�%����u�ނ^��>8s���6CYU���ފE1�UL6��1}��U͠�q�������>��4���B}/\�|�{�]B����]*}zӴg��ҹ/+���Bɝ�̝�}���נ��`H#��A��zd���^� ejA�/^D�.:޷Q�^N�튀 0*��"*��U
��b ���$�EF�fy�P���.��*<;���ZL�/��{G�|#�*V�u�ƛ�6��.Y��=�2�Y������f�例�ͪ����!���s�!�ū�_jy_�d<�D{��u9���Sc�o�Q�Lg�D�)�xfr���%�L�fy����gL7�5��xI��0=9�a�2l���}'LF��j�/IA02��j���n7&+���6n}K������a����|�-f�=G��l%��C����Z�_������ñ
���,m�D�h�XѭYw���J��)�NN��0WQ{�h$^'+�c3I� �x3��6��J�P/�O�Y��F[t7����u����#�w�U�=�J��5�݇�y�5��m�TrWn��@��7��Wju�(����w�;,��<�߻]m���<�A�?�D9��'���r�نMf���j�&��|ԁH�%]�!	l0�YP�hb�ȩtf��f%Y ��C��=v��3FQe�M0���eX�	Դ�a�B��9��D��cv�	�[�x(�YE����ym�K_�>�煙R��V�&�<���o�9Y�S/\�4�F��k����L�����,�1����ڄk���l5X.��A6��n�!�Bp�)�5�D��jp��X7Z��O�~�$u5￢�{e�V&^n��+7>l���z;�F/��Q��y�*n��&s�/3N��8���8s�N"I��dj��/���f�lG��n�,~JDD��#(�g'�'oъJ7Ɩ���fUȉ��W�l)��ۙ.�"�/
gMh�R)u&�n�I^.DNm�e}s�Re:M�����m$g���}<�[�(��ib@[�x���?���-�������r�6Y�Q��p�l������?GV��((�c������Y���,�cϗ�p��Y�I�؈i��z�8O��[V�.ʼ"�$�'��c���$�s6�d��	�U�'$��CH�x}�)�J�\��\����:��dd�S���5h�)�³�������Jk�r3�V�����dӍ�����G��\����"c{|W#�=q�0~�8q3�JQ֔WB�[�����(:�E��|�\�z'»�}i�����˵��-�d�����ȡW����}�^[1��^�p�� �(%��^�a�#�K����>J"�!��\�!�6�..|5��<����bkyh�>1d1'�Mʧ��Q{ģ�N�#UN>ʜp�YvW�]�Y��M���=��PEsV��j?dt&�\�WZ����8�lꑦa]�۟_t���|��� ����ժrU Οv��U5�q2��<�Xu������;�%�9=}��ЙD"gK�����+�<x�㣫w�%��l��w8�ђM�d>�zy1V�b�1�B�a�2K�f�f���³�;������79���o���%�Gd ��P��g7~'<�=�Fi&.=0�-�i���|����(����:��=�K�aJ>��l��wL��)�p����39��eY��<�G�۽sZ���B���t
��`]1��ޗ�.Q�h(Yxx�%~����pke���n嚹.XAڎ5�h���9;�B VJ弍l�z�\�� 4��+qAf��a"��{B�p
�{�;]7�7��2��ˆ�*������"t�A�=XƷ@��[>�%,��p�[�5�&%�� ^�&��9�,V`1kn|��lE����\��n�A���s����\uS��<0�Zg����R���$\Ҽ#��ɊSњ�#��N�A���p������R��J �'`BG�pV���	��l�������?[�S@j��<����-��+�}ɓ��βJ��h�[�cω+D����#�虵5�wa�U!���F�~��u,�3���0~p6OZ��~����n˹��ș���y1�q{��J�Y��CrS�<�1�CX<�j�ب�3bO�7l�3� �
-�T��ԧS�6�.�R$ʖhug�'�	���X8&���?�i)�+s1yZ{���J���2�z�9��,�lX��&>q>��e�7G��;��uH�Ж��p��Ӹ������۳"�F��2se�u+Kq��fx�먫��S��+�h$.�;f�p�fǓ��C�{C}M��~@��*���9}�b�`É#�u�W��"���:t�k�j��ьyQ���ȹ�2?�m��,w`q�l�Y��!��?�#� �|��^=�=(�6!y�OY�H�z0�����a$�
On	~�VT��`��x�XW_�?O@���aL�B�}W>XxQ�}�:K1k�DR9z��U7M�p���������΂`x�X�o���*K��d���;��s�[>�k�y�w�D�u�]g|_�j���Jei��>��IC��U=Z���竽�S2�!״���Q���e��(�\*��* M�[�xgW����Q��̢�� f�ʅ5������Ù��!e����a�޸�,C�oDK��|j��w��s�n\���N�l��s�)"�JZ�t�'��9���fH��IOE�X?jJ��:g�~�K�*7���f�x@�6�d/��=��pZ����v�f��9�[k
��$��:�K?)��F�P+��I��i����^o�����Ə2!�f�Q�F蒵8�Xu~P�R�{N�%~$
��2���ߪ3b��W)�V�բGiYZyj�5�����rLpv��J����Y��
p�*@�[�ں������D���.d��M<U�q��r�C�,Vo���	�h�{�0��tD�g�j�ґ�Q�FL�i/5�4I&d�����Td���	ObO��ب���R>�� �_TM�h����cT�7�%��k=!�bGE�m����	[7q��@i�O����7������i6� �wM�V�rTW��|X�h��b����?�_m�*�<	_�t���d0��P?����p<�������g��:��r���:9���b�I�O8ɾy�aV�$_��d��N2�V7�n���B�b�L�/���4k��W�Ī�ˆ�2Ú�_�ֿ���Y�?��5��߄�;b�Vݳ�O���r���0Lo�b���e
>Ɨl�m�ڊg6��o<5������HG�N�����jׄ"N����~&����@���J��^�'��S��R�c �����V��rݻ܊��������n��Q�����׺�� �_h��Oځ�j�Hk3m���ݝ�~��v�|���}GTu�6=�����9f�i����G��}N�_�ן]�7�1+l��#���(Yw�2�g�m��!T��!I�iӗy��$5�mI��d,�BgR��-�P

NH Z���Y8j�j�+!̉M�����@���ߩ����)2a䦘��a���넇Z$E����ۅ�i�)��F� >�Q6��W����6����s?I���9��)�� ]�Sg���9�8���N*�~^"R��ɢ�3�9��Lb@˂��W!����/��l��k�;���kd3�bЛ���ҁ�U�&��{wĚ���>')���Sh)��e����Ca���
�n,]��y"��M��Y��h�F����y�֊~��iͧf֛�}"A���z"��K(�/0�x[��|�O�mT�F��!]�{b��eI���cd3K�ɞ��M9n�L���mwjiY+Ց����c@�n^:ِ:.�6�lf�w���Z�~�����l&k\ <��5Oi,�r�M����/J�r/��*�q��ڳ�=%Pxp,{#�!��h�2q,5O�w?�B:6��c�o)\�٨w�F�uo��Ӻ��=H�gO=i��j5����5�u	\h��+�C4ܣ��2��0����*>ߘ�*.���Q��)��/&	��X �Q�����@B�ήa:[��Vu��P�jF��[d���������g�8�7+�~a+-]��a9��~�.}[��3�4)�><w~+t���7� ��/D�M' �h���@�L����<-H�)���<DwF��q�O��'"�����ˎ��*i�p�Q	�hE�}�<M�Q̓:����G��S��@#�2�,i����l�I'��,�w�b_��Y�YBĠ�ķ
�L/
 z5�gPG��u�*h���z:�<��~��[�b8�G"c6���V�Q=��� ���A�O�9��G��7�E��рe������@U�x0T��棹dKj�R�Z��M,G/Aߵ�ښ	�_	�D|���4Z
d^hc��j�h�Z���x�`J��� #�ӳ�/^2�Z�`	�?�7_3��������M��TM��5���Y�^B�+F\M�7o�^���;�Ȩ�wi%�5��x|�M�Y����:
"����9��d�z����i���:�Z���6O�� ��۬
�=�ZOS��ƹ�(�����*�b���@ښ��	�{�6!��B(v�\\y;KC�k�Fܵ���c�4V�xƴ��(M��I���S���H/�P�S bOw[�fUm@8����T�	dux��9��)L���>����4h���V���\y�v��,��AY0:&�em���@�Vbtb�Q_�����P-VԚ1�5��g�g'���'�I�G�[�Q�O����"�T@D�l2��硶��C԰�D��5D�h�P�D�u��D��]xO���L�"
�~��E4}�wcx�(#U��-�.��ae���X��T�5C�u.]%�L��lÔ�d|�6ց��~噲�,M����5��'PՀ73�½�����3�'(-��㮛٫_��(ݜ�Vv��5oL3S�Y,�96@h5,��r>g�_��p�n�;����?z6/�3繠�U��n�E� ���U�U�Ϡ����"��=/t3�R�@�����h�9R���KR�l����DQ"���mUr��R��bpbre}�zn����}���E�x&��4F{�Z�� ٘ygk����c��`���h?���ɝ��UQ���<"���Cӗ�|c4퐭��R�-���fō^�!#GD;�Sf���Z�HxS�W؈k�[�rsƎth���-ĦlPx�Z5o�¼a�yb�6�� �:L/b}��D#	j@~1V�ݐ�4���Z*�Ydiނv��yY~�r��Eo"B�6�Y��� ��"�t&B�+ �5�;3�u�o@���5���3�A{M�r�������.�>��2�>�x��}��y�tg�Ȑ�������c�$��o��Wm�<+�W`�
��@�ĆTd?WX�x����7t%�vR�~�!�j[�p83v���brVj5�h�����d���gh�.��+�IWř�E}j��3��O�.y����=9nj�GcWTh��n�����p"�;��y"�Z��Pֆfvasv6�������j������dU����q��Y���{)y�H������І҇l����IG��2�(�� ;��ۗ2�E�r���`�=t�R�rC$�#��0�����D?op�+������.4fv�o�IiM���&���(/⭔���mQl6�`��?��uSyL{Ws����J�q�!d�=`����!?��$o6=�g�Ǎ�f4:D�O�.5���W�<<�B:�q��5����;r���-p��d[Q�Y��Ir�tN��� ݀�$e�H
��m��O��6mU$�BB�M���xw^֗�wW���Զ����*�Dd��DK��<񭦧�Ҡ�2�V�h���b@�~��>��^zi�_\d�:a£�oƝh�}�19�9wI-߇19_��T��6ȩ�ZܤԣL�q��Ԕ�EKh=��î�W ���V7.$nC�����t�v�["�o>k�W�,���ݏ�e���J87�'����`�W��|�kIB���Y��A�N�}��L�}`M��w6J��Nt�q>*���!�:ӊ�j(R�!�>Fc�����L�C:�=�#ݩ������gг�z�	���2�k��e!�q��	CDSà�DGU%;LW̿`j��X�r�%�������ƪ�U��Zp�q�~s�Pb�t��+�z�m�`+�¦���^!_���������O�L�� ��N"g��Xt���be���[�Q�u�"�+�����(=�np����12�˿�P[7K^a�#E����`Џu�O� )���Sak�U'����S����?�I�V>��K4���U�I�ş��4(��p���"?�ݸOY��bP%�@��PF�i�^����'�^r��+@�2e��s05�N�|Ca|m���?�~�`\f�&�S�٧an`����'��;�fHq+�SI��ኣ�n2儂=�9� ���7�ڴY��UV�`��-=!�MK��H���揭�7��d(�Dg����^���f�e�O�Jy�R���8�7`\(�),�"R��To�zV�30Ϡ+4�bP�B�%��R��l�a��^QN�]��Iq�e\���B����'�m��-	y�Ou�g�����ױ�)�%�4x���]W��+=�@)��]{%�D�u����!�T�ѲKmC�E�Vs*��Z���l[|�����4a��l�J��QOS�$~���7&k*q����z��З1��T$��bg�����iU�ά�����lsP�����?�O�tK؞�1�#v[[����.�X�r�ܟo��x}
/��T|��b��U�w_Ɠ8�
���C� �8�մZ�C<��N/ʬb���R)"V�?&tO"4<B�U�r}gN��#Z���[RK*h��ۥ~�b�wՆ;D^l�0�
�˲�{K�Γ�-�=\`sK[  V�?�M��	�[u$��ȣ�G��u�I2��t<Ǌ���M%����gƯ� f�]����	3�M�=�$�Ւ ���~�`c�K>�0�-r�"�A�HI�ur��t|d��V���e"� �?u�I������'0xӥú9	��I(RX,�a;nkҲ�����;�c�4�eK�t���	4��j/�4�!A�x,9Ew�5��~S:�� �"�8���f��LSD~��f�����6(;�F�rA��u"іb���ko�x�_Cu�h�0�҅N	K{�{�;�-_*�ה�B��ƌ���աM��E�Q��U�H��6�k�-����r�>nq{�#lUX�#n��c��}e�O���8E��1V�=a�-�<�qF�Xn(��j#Y��� �
\��'xpy5���H������3�>h��GɎf���8.����3Ǎ���;�_>��;�=ԯ�"y��e�U�f�<��/ŏ����Ń4䋃@��eJƦ
|�!������:�j-��廾�� ��S��|-�l���_;ίZy
��Wc}�ɺ`�<Y@PxG�:FS)�\t�2�J+dN~P{=����A{+}q�����ɣ�2|80�V (T-��2�(S�ҩ՟���aqx��_x2YU�L3����Ȅ��V*���2�!lu�k΃�����)��S&�L&~�$��v���_RW�9g(8O7�$�U�VYE�V�ua����-͖+��}}�S
�0��-�����f���hR��)�S=�zy���l�m����W��9�^<�W���ac�b���u��"�#AsV{����� �.������OP�}����,�\�n!�N���n(�0�
��óҌlި��ʕ�P�U9��[�^T���Oաz�3v�
�Ȧ�;��d�,�S��2�.$�Aǒ�'S��uM�f|��.S�<l7z*��G|��q��&�0��D��y:McӨZ�H�3/����h i�J��fF:����8��4��?7�Kw��*߽@�S}�m�Z8T��Dc��T���J�Y�5�pw�%�����)n����=@��+p�$%�3��YTN����xF`y4Yg%�:�F��s
����.��Oe|��N��}q?��%�P��Xv|�JUR3�/��ō�jE��o��!�=����8��T��7H�����ލ����P�MH���_����Uj�J��m�e��'w���;uj�.�G��e��:G9��G�>?����s��6sE�TS���ڛ��J�\������7S�ZC��1��q���d���?��Tq��p,�=����c\=j>�k���>fdԁ�3QF�UεO�B=�c_o螧�ۤDF�#�R<vq�>��������%(��b�
�{�M��ډ=m�p��E��L�L�Q %���yf��6�����6RF�W7�O7�լ$�8����s�q��K��	���πi��O0�1u���{��'�:/�,��/Ȩ�p�D́��I����M������?Ӣ-���ʌ��Z�k8����olwz���M�Y��@A-8B�����oOf��}�ˈ�W������'���r�$���Z:����і.���mLK)1t�9	w#��>��B�:�H�U8[@dMXR���e��<@��U�pCR���]��K�*Ēf������pp�_�qX�'y��>}!v����?�h���#|��?�O�+_�J3%��_�Cdq�,[,�J����ˡ�x���|����H�}�E��_L%��� `���|�}�vv��$�΀��@t���J�v�����D����e�˔��@
��i�IE'C�mb[Is�i�Ԕ$��W:�˪�S9쌯U嫳�E��Kl�B����.�ݶ}p�{R>p�|n�� �e�挈1ju�j=t��tG�!M<��^�6:��ߥB���!e�X�9�?I��q|Z����Gr��
��Z+vо��F�6ŌkX��^�����+X�ۺ,h^J5X�D%N�Cu=1/�co��~���gM�O��/�
���xLfmb��7�)��.
$S�Lب3�����d�n|%X�RIr	���\5
f��/��e2�_�.��(3_���"�j��u������=c-��}�&T p=�]xRc�M�/&���ơ�"��!:)�1�=CT��P��}{le��B����J��{P��n"DE�s�'���qߗl���;)�MB����D{^���^�/O�4��M�E���Еb�|,��ֆr���'�3=y��Rg������������k
����fX;��������Ehx̥��9��(��v�ms�:DG�&������ideCE�{��e�dr���8��+��45p�i���r%2yL
�P59�J��$��"��tv�W�9���	T�l_5QW�wH�a�%�0TZ�Sa������k��7Pa��dC��4[Kڕ�|���+��Uf�I�J��L�QZ=�-�	M0Wd.�-H��r=� ߐ�����!^���B�x}Ă,���!��/%thz��6�g
�q����%����d�B�ܳ�6/��W�;U���(��*�-szj�V�&#�{n�Q���&����ZzIw��$��c����a�A �lX,��E�����GA�Hk[������h��7���rh�0N��>�=�3fB��{X�i-=(a�&��R,��*�];�mր�b���S��1��RP�.���<�C���pue���Y����O�������8�O�%�(�J���1ֽ�q29�)R�����G4�\R��O	.:���u6)��|��݂b�΢{�v�R.&/*��=~��`E���񿐤G��"��c*����g�J�ii<�_︵Wb��>Y\��ʇ��Ͳ�^�Wq��ڥ��ܔ��~%���iO�T�����7��0���=�N<��|y�鸓�:�++~I���<)�=�j�����;�B
���+�r��a��t���0�۴�N[��v��n[D� ��(Q���F�2ip]:2-< 	{֡{(�ҥ���Ո(��;=�@6P�{P �:�t�Ď��X�; ݰ��,�3�����=9q��7)<�2j�4���L�����Rw	�J���̙���&X��cl~QE�&�I�=b�V�F���6����vB����5�_y�����Տ�T��L��uE���j��!^���=�تcZ��D�~���_��CXA�m�!?��ᗁ��[����T!3;D��Y���,��+-VJ��N(XHT`z� �(�����u8���(g%��h��D������N<}�l�e��خZ���B����}'��U��#P>@f����%a�9�;7����'����.�zO<�6W������Y��F+��]�J�VE�J�v���LK�.`��ǫ'�}������2x>�g�'-�c�bt	2=�_�/�G�8'��w��.�~1
�nlr��b�~mKC˸��˅	�{#ɋ����	9���)��ܼ=���M����4�.����u�@��܊�Wq�pq��y�XFC�4�z��
a,�d֠��Uq3��y�	��\G�ӱ�Й�Aȍ����M3q��p?"i���dT��gn�ZI����%�1?�w�����+��n��ᖷ�W��Q;��r^G.�-+e�qvؘ�i�/�"O*ߔ[�E�k��N�Y2�\�V!ت���8�D�+6` �>���;W��I�5i�����>w�lKl_������7�G�}R���m��`�{:Ai��l�
�j��Q,C�Ke[����`� 1��@8�z�v���D ®^G�����ӷQ��=5�V5�����	wx�`�,v�.a�5+��ǉp�D�F�O=�p�O8/�p����5}�}u��pز<Ԇ�X�#� �0��
�o�ױ8�m�R}z|������UdE��%����H)�ͬ��?���f���� ����h� ��F"AO)# t+<���X��Y�H�&�������~F�����|`�Y��s���[�t��"��wR�y8q6m�ST v=u+,�`9=����Uy���G�&���2e�Џ�w\���U-��N�m���t��(�ô�C�7��5�:�.�O���N0�]kMΛ~��u��������:y�9��&�����A�d#YN��	L�vu�����������X�i{��Ͻ^>�Qp���m'��\�����8��:�A_��D	�|���X������Rׂ~)���D,�w|����u�6�0�|����/\�T������[�A�q	)]�Y1C�P��I�����'�}�I=r~��R w:9��$r�`���(����2�pl�RQ��H�����h~���]��/|�R.���.X�ȐMk��`�w'd�d�:����9F�������* �)��%��-U�ZR�i���Q���`jSe\�|ha\M���������n>�*�������y����R�;Q3�V�QԜ�JJX]j6W���S�$v��H-P�7G�@Z8ƾ�x��l���r8ڱ}w�+e�)j��-8��l���o�Q',��������a(�z��a��~xГvNC���v���P3i�j��t<��c�N+����?�z��_�۠��Euv��������e�vFΪ�X�&w��>��T���BNz���T;��>�0��'f��b��[��i2G
4Q�7�@�*鰁nx�V�h�\кd���CS�B� ��j���99g���ћ�8#c�x�YHԄ�Bأ�rN�	����D�cu���'�ۺ]�QҀ ,�&��n��L���"�çF�]6�K��?�ˎ��#���	�@�����3���.(q�`���-�(��kՄ�Z5�n��[�wó(F�n��
X��T�?�ע��:��.S|_s���.ӹ��`�Z�::��9�]��J`�}<��g�m��D�����/������8#hj�D�!����e5�q��|�A�M�%U勎��'Wѧ�[����Wz����|�iH�	Ḟ�.ha�����)#���j%����߭­��C*�ӑ���6��K�8���r$b���N��}��p�̼��z�m��n֑�i
c�"B��+�+�#x~�"g�u�w��LU@�|k�J�Z9�zC/���cuFi7A,���O�Pt|�d��x��8�P�Ӯ�P�ݚ34Ӑn\L@�JAGo�,����2��I�X\�+���cR���M��d���t>km�W�5o��D`)�Ɨ�^J8C肣bSձ���q��m���]��'����ɰt%�J����ʈ�i���ː� /n������6&8�鴠�g�]ٙ���v�kn�A*Ll2��,±кL�94�J+Ϭ�1M�2R
��=��@�̇� �W�Ȳ���9�{��?�Ҹ�s��@	wS���)��۽0[O#��'�J�i��>.�!	D�ߐ����Oo�a�jhT�H^�uA��%C�l���Sf0�ʜ�;ۣ�<��9���1�M�k?�Y���%%����gK���E�Y��9o�&O�P�T��ZZ�3#K��/��e���;Z:9��.��յE���֝�E�p�w���_Kj�s��N��� �${�H,�}hO�L�`(�	޿��w�]NF|� ����������e�Ϳ"���Ɓ���\e��� VS�
�=��f��/�v�H�Ӓ��=z�V{�%X\1E�x �U�f
����U)>������y�"9p�h���)�&If۶vu-����N]�����/y^��~^K��{.]��E������"�F>���o�����?)@:�*W�4g�Ş�¤�2����� �%�w1}�]2N��F���Ukt�#�})�U%���`���c���q3��,L������j" ka�iz�ݦ%����kEd7:E������.�vv	#���ާlǙ-"����� �&�@W~�U�/E�E���!��f��	�n�׊{E�O�_�`�kzQ��+�u����yy��<)�����/�EL�wU�-�-����Ջ��pgR�2���Վ�y��C�%�Tiﶅ��I����[�vsSN��[��{N/�P���e��=/@�
"���bv���D/�C:|�*ԡ�5�I�`\!��{P$T�S��we@�1�W!Ooϻ��(d�^�F��`W�S�[')|\D	��TQ���F/ό)��H���� �i����/��f�:x.�s��<X��a��!Lo���I}8�5�?��[/�J��p��+�X�6A�O<�jjPe�g���)��m)���Rt�:/�O_��t$?�1��wB��߁��̀ɯ�0y ��hٖj��k�O�?�<��2`o���%�$p�{&��#;$�����mg,=����6�OI�����ɝ ��ުY�~C/���_\�'p�J���LF|��d,�)�\��Ŕ-����^ŉ/>�#q����5����|��i?�,An�0�������m̿Hѧ����1�2+:h�8!X;)92�6���8T��k�y�|�9��UoW��%�����@�Fx#�s�tUN¿<���J{՘\��ǟH5�k�`�0%�E$��#��N-�-�*���Ae�;x�|�]%|�0G��Ա���Pq馄6NP���;Y��p�S�xB���y�E.��������^n&����pO�E�٩:�{&��g��|o�=zU'����R��88�D|����lj$�<�!���z����znT�aeP��u*�)-ߤ^:����uo�i����نk�EQ��τһ.]�ӌtP=���u��Gm$��~'�/���{��N��Hg�����> ��^x:�|>��p�_)4*<b���ݚ=:��n����;��@�)ڍz�����vNO�{_G� #�B�a��]�8q �T������c'K0��}	Wi��^��۵����O?+�o�\��\�:D�ݓ�"*d��b$Q�m�ԩY��/�\tF����i��������LVc=�y�Kjɤِn���'��]�cÂ@~�P\P/��RӾ��9[��N�qwft�!��y�P����ǫp{��u CV�pݹ���V��hP,�3Jȡ:c�e��௙�ܮ"�lT�S����y�ҟ^Tm	��
T	/���' zk�F��w`2��Q;��6����=�Z���V_c3z�x�g�u��sh�Lb,<2H��e�K�Տ<���#�N��>��V5��&'�i9��6�Puo����0]��Iy��w��_���9��m����y![�>z���LT5d��r��О��B�M��Й�0�7�ӕ��<vע`h�p��|�كmny�������>�'�مqe�S�	�+�-r�ɐ)'�u���$��d|��7��T�<?!^���|��X��ˁ�zlgYJl��Y���r�_*:�unчyL3O��<�V��"֪D�u���A�S�A���1�tS]Vq�mVm*Q� ��JV�aJP�3��ȝ\Ֆ�U�"������� ���aH(�a��1�7|��PY���z��X_sl�X�����{ނ&�3�i��Ƣ#�d�4Mw-�"�E���83}�H'ɦ��!:�2|�̈́[R��_7X��\� ���OSA+$�D�$G �B��B�N�!���A��Y����3:�
neJE��mH����Ϊ`��@���ґ�t���\��	�م�Ƌ�_]�����+��DI�
�l��>�kz����?�$���<҃V��	B����'6�[�}�"�����j��o�e���5����(��/'|�w�[R]<�ʬk�4���A���X��~f��ț�Yw����ݔ�C[���6�6O��5�n��1���$~�f���T ����#��@��\8@�Uj�~�V�	о��-�o_&[��l_2|��:w��[���|�%�m�(�t�o�E����^Z���U���ޅ�����x�ҩ�T�汗�C�̊�t��:��Q߸��♓:�l��ǰ�]����*#��n²�z�}$O	�[]2�İ�Oph����F��ui$���#*�;ne!�=�Pt}�&lJ��M�'Q��U�/���Q��V�aB
s4LӾR�c��6IsT�Gx�X���������^]YQ���0��v��Ҝ��=��d>�U��y�X��A�$̱v 8��������i��_����_Z�}#^�܅�$eJ e���؎l���ntKR4�꘿�Ɓq��\wj�P�'iئA��"�#�Q4�NoY!�y@��f���b7
k� e��ڈ�:�ö�V~��#[�H��)ƹ���k�e$��H�]"!*� B�6Y>��H�쟭��QE�.{��a�3r*`H�{��Q�XS� |�.8�*
��3�h�E�pI���s��_C�`1�I�����):M�a���"��fb���j7���a)�	s)�)�u�: �pE��ѹ��q[��)�lh)�NI���֙5��5Ϳ��(���=#m<�H
���0���\��F>�.�X?t�E��$����O��!��Y�{�z�t�z88�5�Av�x	m|q�����.�=��ȶg뺥[�Й9�w�&�{�p��M5l�������HT*�ݪ�$�����C2�\����q�2�J�������9L���5���RƺS��(�23QW*�L�:@YR%��7u��Y��I�Q,��O��##e�����AT{q(�����m^7S=F�a���߱)x3��wŇQ�"���^|��R��`m��p�K���k�l�^h�X)�P��t�P��de��)wfC=��y���#����[(k0vXH�~An�R�|޶rF-�ު_��/��j�#�3�}�O�kv��Zug�5�J�0^Q>�ն��b�Go��0���C�ΖYn�{fh��L7n� ߲�Fw?xm��e�M���&��(�+w��|�hV��?'�^iE�3�}�w�ќv�Ai{�b���Ee�s�aBe�+V���4�"Z��*��g$Lj`�1�Z�\���罸���!�͜�906��x���w�/Oߵ�B�H N8rD�SxY�
,�:���K��#���I4YT�;�wR�|����7�h,�m:����A�z���e�����Uo��8�?l�o�ُ�GR��N����z�Z͕1�3�}��o�L�B�o�l3X��Q��Z�Y�pTZ�)���H&'!��+QX�C�����@#B��{��>?1~T��
8}p�':�[���y�k��`*����%=�l��U�r-F�������w�pt�.��V���Y~���{i$.S.��_��$Z�W.ɚ�5~�F�+
�u9O��Q�X����cLj�pB�g��9��lxxc����̠j U�}��n�{�A=4�t�S@��9�G#K�]"ϱh�b)�-�i?He�/I��P�n��g�.+���h~�k�ɝO�t�
K"�ż����"�Σ5v�w�;W��s�#	�j�A��C3a��TG8n����}
���z5���z;��׭�h�R�"z�
�q�dF�ܘ��M�,h��k�^T8�D�E�8S��eK�qܲW��l@C�{T���#�H�o�����O�����V�B�p�rc&JJ@�9��ԭ�_
&�"~���Sn;���Mzw��n)K��d�Qq?G�ƛ��1��ELo����Cz"m���#R�g���:i+�3�Y��2�APE��|n�uV�ӏ�8c� ��C��&���Dq�Z��LoV^�E���N �=`�j��-ʿy�Q4T���(��C�d7*��$Y��,0~��fʬW�@~�+U�f��MI�R�g�ۭ���7�������E�����Gj��քlx� Wҷ~��#_�nV��Q���ؖfM0��nG�i��:�/H_���o�ojc���*%F��t�7u,Zz�A~AW+-�t7tN���j)�4���q�����^ʟ���-0�T�,�Z��<(�H%��Ws�?��+FN��´�����R�5g�o��)��^�p����C��d%�w%��P���CH�ϰ瞭_�/3?�`[�����B����l�$
:{@x�� �:�UR&�����q�6s}��L)J���0ח�_�~���83#��1�*peU����h����N���5��dv���&^U����z����Q�6��+�L��k��	�+������~�f-�0a�_�H��//9���j$�t,�Q�(n�)��&��1�1!&n�\v�	0�F����z��Q6AF���u�~ݚ�}�Fl"�Eiї�Reg�f3j���z7cc��iއ�ׇUۢL�4���HIC�*��.W��9��!�c_Q0��J�e<^�&Ȣ20Q��~+�1�n(+Ķ��=З��9�M�� ��`�j�H�&�9@Qa�^��x����R#Wђ=�����>=�޻�a s�_pzS}Z���}�fO�~I�xĸ-�+UL��Tl�E��;�*V�[q 32 ���= =ų�s��/|]�����ꢶ�+��yfY�{�+Q�$\C8��]S_�t�d�Qű=m̐�:�-���2��r]���] gs�P��[�tx~�wk���t�Į���o��.����K�HR�����D���dY�3 ���g���$���S�s^�}Dx�ԲF�a���x�J��5���BUmuIÈ�L_�T�}���å�����7j>$�M�uU�Z֮O_DP���h̲�S�/:`	�T���A3�9�4��`�!l���9��A�'7�Sv��'τS<�bs�Z���x��G�'�𤥘��#�:�G�����8[	&��=�p.�խN>ރ)6��{%X�:<Z��{
�ZY�?��E2�ٴy"�
��q%��߸������7�I�T�ia��%]}out��PTJ��l(=�b��ب,��N ���s����YP��Ԏ�t(�*��^�?Ѯ<M�s���#ס�b��0U�������90n/(7���y��P�x���q����ϗ�EǹU��y]������Z�d��q����ic���[d��y�۝xnx�aR:|i A��VVc{�6��\���\��\R�'�#�8�u^�l-��s�Hd��X/�)�=_�p~�l�k-�_�"���݃�B�1&�G�Z��/��o=n��F�>���]~)a���+<� �ab3��^Vt�[{� ��YwC�M��m�V; �侴�������|̅�\�5�_�_�,���S��ɧ��=8��N��b�ʫ�%�dw�C`�PS	ƒ�����K2(3-{1�suA��cj�,LT��,�ay�n�}W��NtG��!¸˂65T�=ƢN~w�5���,�t�ԟ�.J3�������_6����u
�[��J����3��}z�i�=��u-$}�5�В�\�B�c>�%m���;���mθ��C��紦�&9j$}�Ԋm�r��l�u�<��a��R]���d�3H���5�_K�@l�2����}[*@F���?�ET��MV���@^�XB�<�Sg���(*���U;�uT����؂**&���k��2�ғ�_����I�שEF''IGU���{���c��х�;�?!��W�"��ZցJ���}2�뗦&u�k��߬��p~�g�0;��X-��٫I`�)㨛g̴P��kEd�

��ǙG1���)n�8��G ��aAd��9��杖���5%��]]��VVă˧��:�e�C/��q#�*������\�nO ճ��+��<�w�b��B���>��{����;j~��L|P#��[�vbT��w�������R��;8�?&7Ҳ�D%M�a������L&�[�����;�P_f��/����Md���h/��wxSr�U��ݕE���~�*l<�a�	�!��^"#t����W��!�N�������w-)�2��$![��
ds�|�f;��61f�3}6����j�O�aQ,�0�Xo�/�r�^�/h�j�	����f��A�29.�~����.P�6��4�!K|�a��)������Y	E�	�P.��6�<�2"�=|��h�~��5]�W��#9?�uu#�tk"{Wm�Z;~�W�m¼�e����]�;u��Q����b����Z�������a���5o������if ��p�!����7h�.��@�"�SNIYe`��B��nizUbR������]�q5�>��S��|9�:HJ�@�]�"�R�,ްF{$8r��F|�^4�ͩLs�V��YM_��Ibp�l����[�@t��`Z���o����r��i"��.�6LB�Źb���e��0�D:�Z�U�R�Ly�m�[,#�Px��Y���.�;]�|���F��/T�%]���v�2����/���ǻ�4�mz�2�:�4���/#��$W:&ğx֠"4,=m����T�}R��i/�` ��.[����C���W�Q!ҞCL��%�b�Ȏ4�u]��A�T���S���B冼��
�`�:q9s�1����0��%���e@�q��f��-�Af{��p�ߐE}����N]&�u�M*0��~�W<Ⱦ��%��wm�!�Y\I��p�\����}]{�Ӵ}*\�Р�:�C@�&Z2�=��
�Bb&gC�^Y}�U�𽃏���z�{a�3i�.v�M.R�֬�RVꑣe�+Xw�P>�����a��A��ԾD��qTl�W.L�k�E�]f}د��UvD������@C��54���O(laī�&0�9�՝�ӍO&�������;6�^�����=�lFy����)�D���._O?�(�d6�}�M6n
_�za���LB�����D_��9�r"Rm��IbO�p�:�jS��M���B��^w<hs̢iXh�/�%��I�O��j���
q>����z��!�-�d�6�Ii���������2���{����Y���-��9��q�Sɖ�靼]����E���L>l���%>��>'�j�n�-����K������ڍ�L8m%�0���T�ƣ��q�O�T�B��{/�a��R�OX�B��_���wT�=)����຋Vk�Jfr ��O�ݹ�]2� �21�u���˨�ѩ���*#���8���#x�-����߾Ya��|qm3������c�}T�[ChgET�������k�����-�R_wc����8��� ~t+�\�Y!bi0����3��p	'o���3�:�(��]|��6ᳯ�6�_�܇�0󳮢bڈ���(oO�l�Qʪ��D��?Q}ނ�Ő��ý��u�b��x�������Q&9A�|���	�\������7��uN��jr�H�zg�