-- (C) 2001-2016 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
scAM/69riSUUhLCtsNDhTPsXFH9KCV2f/YfwMXDC37lrpLHsw2PHP0YxKA8Zh0XkQiHboMEUkyKQ
vxMLaAUu7XnvUctLHqjR19h3qD+pXDp5v9uIx4QwsMK7iZLkGgDJJ6QjC4d33sLK6PAc/PuidSPC
n/CQ3s9cxRmANiD6qCuSHtrZs6fSvJUvMg16p26wKurC60hXCjXN2QjCFOc9w8ztJL2i6hiuEk14
GhHQMmgysQMPkPtLndEZmcPLLmeG78VHNlzbI1s//S0ZdjBwvsp1dmfnR6xtv6dCkysghFOAq4z+
0/cU8P49Yek22cutfIds23P058cre84+TJg70Q==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 6176)
`protect data_block
HcJUay9zEa6L9mOobXJsvT6aKeditTdzFHsHpczWQFV4dassUa/DmhfkDinf0f2+1r3m6O88shAL
mASZLITE03mBr5lanEMhyMlljnHYJA6VasXDznnuztZZppu9XXgBX+HkjZL/eovZLKfM1VP5TscZ
yg2fWWr6JOmk8/w4lpIKDEYpoPfYpLyFhTFddMtlyvFYsul9tsD4w+0ma8U7yCqtbjxw0hZr67E4
k57usR52f8So7MU30Swott0an4n+Bmstn6flQqiXO0F3KycUJLmL+zMjmI4/UU92CqmkGKaqpnC2
igH7F/3sR8Mxi2Ug/h8v04MwGFrFNplg3j2vGcapJQrpE6M3sGjEVqrifBvKpysFzR4ulRMo7IKV
m6BvKXJ7/hiT9/AcbVpavtxuElg5UdKcXExRDK3k4oFi6OAW2HiRdRfjmQLgmHo38GA/YyPz3LAx
ljq3L/D3h5w86ggqgKrXrFTgkTsqWxaAGzcFkwp3+W0gvQ7IH2qT3bxpVApEIevErxx3MV8Eey25
NGSDRMSXdt5QR1lqYdmnIgNJ5AKyFv2soppu53G14iy0u7vrapYyQcXLQRuFEPmSWEGmTZ7q6nuv
Ny/Ogo7AqmP7MnZgndHXKS9nUjZaQfWPT/VMgXgMM8CGVnInidOYcLJyvdS/xHUEftQqkUJ4sPbX
7T2qpv+sNtxO/CPEAx92ajXDUrZ2xfL+9KibMSoOuu+OMtSlI9kKI/DfZU1+gTkgZW3PeR6vpT3E
SCyzF+RusAH1TJnC9YmAnntVEjqTSIiMPPpil+o3WZ2+dWD3FQ5rjIcjL94la4qxfQugttTanjkW
zOQ5UeMVDr9pbvt0CcKDBB5umaD0P5jtlGyh1hrViPUIUBSRl75Dn+i/PtFEXUBii54kCkk8ODTT
t4bh40E5tzWT7Jh/L3y/iwjADRErP3DnnhljTPc5g5K6fjyEL4BHcl9zrxsJoQMAeVlJXQfvjAN7
2T1yd8ZqpJNJsMwSJ0O9O2MtUi/ctlxkKOClIBqCEijMy4PNCIxU+LXpmm9GtpwSpg3w2X5znQ9C
PtR6EhwMQU1AEJoWZDrhvYgfaE5iriw692CN/FOa3kNSB412f5Y5fp06A2wPitFNONedGOBjHHux
LSFRCLO0kE5Btroa/ReWkT2LrFNPncwxSOK7oxecFcfACxMf8yZSrau/PlsFgGzZxOCaE2m2PZjQ
FhvAPDYSkMUgdZE4XVsHW6mpqEx8JxQqqejtAgtaMrh6eO1ryvt22rQ0XuZwYazCBGgPcZGmzG69
AQoPfNxA21G8djSzaM6levO3+3tP/09pmEJmvGL3z4qtp3jQSnwYYc8+FJB8U5XW52aWXphtLQZ9
39iGitGf1GBuV0RN+s44LS6f0X6BMvN2kJoc+WP19Az+qgoW44WtlZBeD/nPman7HWU0sK6N68SY
VKlKFPu5OyN2Jg9hsWhiMegaveJPkOuchpF2a9mx8YITUyBGcg2pIDgyouVKP5vHUO0I04f1Em/j
fGPIRAZEznvCdniMxhuwuAS2g8T600JrVlGqhh4Cr/WNM+91I/eduAPGSsjYCcjRjJuk0ENtsgcQ
UEStSrl46Nlrm5yjgXQEx7Vcs//zE1/e4fdqATnAcasrv4rUZZz+fUUm5Yw7rpYJjphTs7Q46MiQ
FizH5ccP8RRntwggzOr6nxUHVwU5Mw8f2mZKi5ZhuijbhPkRSUUh73kSHbuQUvba1C9c8LcOHMae
r+ayKxRg1iuQH+fJNAZe06GhKOLW4z8WiFFIOIOOYvthzYfzL+lyOgcfpRk2szbPZDgewc3hFua8
1iOzglBl1uNYfu0yQuoVNjQnDeDs4P26gdpt4vawJv8GQkQG2+lB9CIwhAzqoyqZkum0GDKb9d2o
QX+vNAXlGEQqeppmZvnNXVJXm1H18AclsPXZCE2pODx7XUaQfLq+3xDXI8Ewa/AbU9lsJJT02c31
kVe2GU5vAGfFsrKjt8sdosRNyIVAOUou7HN50+h4JIXvRyG0gYYA81j2sIGqrE4H48jJ8+pZXRt6
aOFrD/iy8BnADvoffZiltGV6033r9yPGGDlHSni5z4SBYOnNgRW/CkqqIMOnOripufxWaSWGljmQ
s4A7kevZ1/tgPEwW1/f523JJngv49+ZUyOY6oGIs+MlT2GUGVYiuX8beQvzJyc2kvaEkQb6E5bQC
sQih5FBspFWoimPHtDuEu0ngXINgD37ytO7RFI21goCHSHqa6QbGG3rofEZKk4UwgKHsRMyOxYpp
LU7ISJioHiZqzjnV8VZE/TowsxqcSCgYdcR6OjOuOpwQBWvbmBHiAxzQPtKuongslqU3R2ECV3/M
wuf1TAUczAcWLOLOp0pvpszh7lBZq7qRB5/rJZKdNm0CrPV6keOkxUljqFPtqDaJiQkxpKz286u5
0Q9OqAGcGo3sY1NVhNJBXXI0jr2Kc7TIGS/4W674Djp9hHiufzh/PBrH5t5wh7HeUdzyxEyliZlj
bbvgooH95l/1cvBc0EmXogwyUs6DO25Ogyz1KZfs0r1dtyAQjIMdG/0QiG2hpaCwvt+BnAgtvtIC
F6iT4ZQX3A34DMwE7aHwbr0y2X19pIp1dBmIHJaE2PIGnd5YAOk3i7k/jWA+wNCsyuToLaXsGI8v
S7iPKX53R/V7dB2FQH7Zs9Gt+9DBd9RRPvNcPU7CJklKPyy0sWLEdg7juCSq48rFErbxGHHKLjyk
v5NeQYTXfw/r1Y7oqIcQor+QGNUeDdSJ4EwHtv68AdNf8KM/vsPwz2/skj5C0+ACkW/PwsjzS+MN
rTKvqQIkaJcAXn9HOAFge/WG9TUYfEdZ+ZNZdxf0m06nFkCr5FZCgpVVHUk8UzmJ7cjgFWl7Z6UV
tepwHEN5HzwOW12IfcFgf6JJl17vywxKFJQBQb+JSQQo7W/k+LUikl+S2Lis1ntkWkz0O58zWRl6
6M80CvfhMb3/cUTC/OtiovJxY4/OfLej9TbJyzgmorP+PxR18hMXc0QsQbKNSNQEdd6lye/XHzae
2B5fo7d5bEPu0vvvJ7kYCqZn7yZYyIC+8iCh7XHfy8EhN1KWVHrLKWfkG0d1QzonI5aEQj+wrUqn
xEi1mvSWwYM9ZiKKvLVvME6/q4d7XlF5X6aAhA06KeXSJw4ldJ1i5jVeQ5Pl3IJfV5u6sD/AZKTz
PDa9YPr0mOWcUz2kCd1ByRGoxebJy/JG6NWphqU8nWFWh5mjp+okiVDGd8QZzfFkZvA0yBi6YT5s
y3IqKpbStNHV2A/kDVT0aiFeXIObT1RGfLmOnrOMrdVg1epBhLm5VtJL0wYFHr/ndMOq7dWP7niY
btXgEfOyqqMyhAX34CZbgnMWpCvVv1nkg5x0umSnz7sfcQ/boRNk0lGN7CFTZVKxwGseTzq7d2zC
ShZkJPzGgjJ9b2FqEoLJDBZ5PKK8mNjhVISRlrbZknVsiVJCS1DcoTu5KMHxxe9Mdfsok2orqu5V
x8r9CLQPN+MXm5qXmaXeqvf/g+5JIZuKx2yE8h81ZglgqsclCkkM43PyyvcWVS0thj5yvC/ijT4O
cm5oOR+X8EwnkeWbXeN8k+O2XNzGB7zvBw179fJ8/ZLgmDMGOM5sPyicRSbsts8RsGYNt/+br0uz
8fa+f1V1QQeX6oMKCp+DMaUWaHmq67S2s+CbGc1CJFSEFXd+DLkMePKiMcMUc8tO0ZJU9RmhuTL0
oWuQPYNJstV8a8Rhs9fH65mhomV3Uonnv566V86xLimo5M97gwy/cZvPMqcOJJUtdmwp4qh3qvc3
lz6Cs/eTh1gFGCLE6LNiIslPNXVOMiU/XRuwu4FKViavOaPUg4TPQHiLYxVUVhxIj9n+EvigBS5X
tQCH72Tgc5Z1+Nw2wS0P9RnQOGqlMxWxrM9a0dn5Kcw2074RuPuNIvz0EB2cUEBcIU9uFVnKDBpd
kXcBhHtKRqp8yFiU6fPkpcOGBlzvlYBmUTa/i6yWvRi/9hpgUvLYuKDiy0nAP2V/0sFBRK26aHfp
5JtE3B+VkgeJ8jmsrs+O/CnU5ESX1WalXO2Qn4isYhS8aMqETVriVR/xfj88xE1SIenqNpJ/hIpp
/NmXazO7J5pavRm0wqABDR5Y/DlIn0mX2PkTZSXiUXEUCDo/XGQTpipUPRmUqJfXOZym8XGR4QZv
PmHzeQSeJHwS04C8D6mqClK9CoBpfTgU5Gq0y7/5U9uWtZ5YQr/MRkmIi4PX2TAueedsb/9EQtoq
NpMO16VNutZGT3H+aingos2bGrbylUBuNagXpcDUBYQalT6157cyK3n+J1ey38JKJZZSghkYfyCK
8tfGyGkRKjYywktQCeERUgVqpa45WQZ/Fc1GWMn6DJNnbD7N04BzfKm06xKB2qK39w4deORpkiqV
sBJEBIcl39W6gqD/whgrEIXDcNGm82XXRYJV9qJlTqW64YLteN87fuJSMTUQHB2GarTfxDxh6U4T
z4xNAhX56dBbN5+9DaXcqPPIAPuo5vO7URkZE4xFR8pSKelqF6y740pX2E5XLuis6iT6+JwVDgII
yvc+xh8I7F28+PEdUDximYvsKHybRxMYMxQsa3juroPlwsONZRQwX7LBqKecSSg9HIk2kUgBYa0e
vi3mPdg8MGF6SQ78Tw7QP0McyUgyy9TeP0sfzohXVM0G0pgW/AZ7ORZv9anAJk/dC8KWe+ZFpGRt
gJrQts5SynjzupxFAMcxWjZPB/0B4uUr7+ketUp5vNA6bkWL6uS2Ksy39LEXRSXVqwRKGh7O9js9
zT401TnZNDi80VRu8NJ16iBd5ZG/zRul46riBGrsSNFJTlMRYmtB39DpOI2BenP9tuoelSC+hhUp
L+78s8XRQxbKxqiOiCY9xVSxnEMYKLBb+J4AJyDS88ldLeYcu6IJTugLN3Khed1NLv+RIEHJywx2
JQmSgin7366f1P39brQ1OHIL84f5XBaFE0s7l7aBmWk2Y2kpZK8RgKgUIWl12WgT6yncr0HGK7Uf
y3Wz5HNvpFqw1BnFgM3eFMQ7ZLVNp3o6C9nxgj2KhJDRG5j631HOXBJOwQUC/eTuOwDBi3/YGrMN
oKRP6N48yFgyPsLcXfSD51blfePU0yaX7fAnQSguXF6x2f4aqDDl239QA7mrzTdzZbpYy012p76x
PUyi91NPRBuQ+tjFyZcfUOZXAa+D4baZb2Wi1L4HKY0o1pr5KbQoHOIYFG0iSitgKPVDg6ek53G2
8HpcKVXQ2mU2yPK3Ph/71T0xNWdbc9rk1ILy08ph5JImuziUenp4YG3yf4P+HXn8V2O6HgpD4noO
1mdPz1sHTTFdv+UOn8T/07bfPn7a933kyzIOAughCC1ZS1aJF3HZI+tWvjVG9D43Nen71lM3p8wV
J0WtMfpp/S0U26/nG96TKpdS2vpbn5YckEgFKUOdvbWfgPS4zlq1zQhHyGHrCgiokKFsLkWCBXqE
RzqfSsMzf/J0XQNFpzZLmuLGceiVkgnzR7s7SdXeF9yYVeLzvXnPbmQeALA4XzNoPM/9a6cUa6zN
rLCXoHcWJQBlwUxnJxqbItKe41u8TnFuAEJsh7lBRBrwpRaCmHxdRC8AjO2mtCwHvzeRBrYPRB1s
TQjRbBPOe72Ryq6I6TOp6FD35Vn1uYZbtmr+OiB/h/W0ZHo/w8Xg4SVEI/+mfQlidOENIbWv38iT
ZSjPF3ZWZhKEhu6fl0Jqld+Z/H1FAi9cu3/pvnntRlTFR/380dQOjOWe3ISmh2Jjaeav/MHjk27O
J4nkGMbl7ZVL5IluF6OObMROe6hmPLJssy355KWW8bqCIaQqrLQfxMHsvTynay4PtUxJHi2/IMNw
ikqR9Q6ThJx13D45Sj4gVanR9hw4cwPJu6jvfcXuI0/D7C85alLKiiRIUI1V3LorBNpfvQyWkdcD
6svIG2wbE6C2hg8QugYFOqzTaQ0HDCx1/t83FW6f74XqeUh97QwE9aRDV5kGLZ/9IU9FLpjXNxcr
xHRf47fyBOYydz3zefLqSqQn4tEGX+IxVRQCWTp/7yOxfb12qypStXm4Q7KltdA67gdXvVKftlRY
/zztbGCPWP63xWa5H5QXfEpSPxYOBlr2yarUOG9uV5JFzCMI+9TSoRImJTpSGmMGzq4KAE3DGEEX
/wGYelFlQrF5N71J13W+Gw3z6kWhPZMNoJjE9vvKL5vno6OHHIgrnEoezMBYDWMdfoNXtCmirY5M
K/+wGd//BhqYttfdo8Ilz+GVZf7YdH/1OlU8qW3CrVbH5IAbgjsxjKeaBzzvZalZ9RCIFoiR7YOO
uGQIk+xbZNFpe/Sb+bUt2K18J5m5qoiyziqZIsN2lNQPWj+XjkboShDhBqVI19WyOvfGU8znaL7q
n4CpRQ0fPgykreV9XGqK9jGF9mw73sOS1CWHGvr+nYKqQoL2YlFRZwZPYe2norHVjOITwwSAKnT6
Yu1LZyTtkALDFZ2J39FCYr8Vp+Od4ENFjOmjlIwU8c84oXBd7G2t+Z4AIFzDz0eEsjgf5xtDc9IV
MC92gM3k+T+q75y3skzGQtZLSGo68R0ERtxmG/PQ+pF4uzrqX0Z6Ar+ggWlqqvA4Jv36ZZXhysLQ
RNsiX6Z7Qf0kMcZkPgicUjKvCDTXfMBRL134kVUgVuLnpG9QpVwxfUiBkm4z2EYfp/9gMeYzZHHU
KQnXM9OIi8fCNwKToccKYtXLKVBEuInnpiEFfiWg2h7r6Vaju8Qu9p4nYl6j1jBWOuI5sLrtc/qK
uo4nexkD5UFrzwZ0YaKHoORAmvqutFsdLyF+CCVEKMrfKGXkH3E5WdqRu4UgT1g8/8toXnH93W1K
OdRcdVb9AqTObys9HaK/X6OBi2MMW+jin85nz9+KSDlM1Jdu9UYplBv2T7bv9a+1mblM617I0ZQ4
n5T894SwWqbblQcETr8I1nzx7v0nwrH9gbCo+FWYlWbFtLxxKA21RPW7y2Nd3s/sGPWXOf1D6kNJ
NsqZOqCIq2z8P7bkEKG71vwv1BpTZTUi6Y12yZA/83NmInYPFMlRh3scwwiVopNN9mNwy1zGFX0p
aTbK8Jvu7V/dIthwJuCMLTFu0pJit2h1ODNR6IDMb0wUeeefhNT0/UiOY1u+hnsY7TnrfkEwAKFm
18nLq9bd/hyZ1lwZzqGkkmMe7tgaGKxTuWmV3LSUGt1FB+dsoOHZqaKMAyyzFyctDVnkGI47/dy2
j8XHHmrCQX9o5oMsyC12r6fBol5JMAPY3p5BituWUDUakmPk8D+NoIS1a4TIL+djIrd2eVlCTz22
zu6qDtZjmF4usZSrMSWMwSE/V5qpXWLD+7xbEBBxtQzfMN7AlYuGvAukFKzZoGE437GxtcKP8rNf
2n+i9NkNOlPMaKN+9/mWs+6vBaR5GqZuiO2yity5IsR6kGsncGGEhRlFr3Po84YbeL8LUxEEpdFG
Jcq2h7QmylCqgAiD4nB2Ur+MDB0E30BeN2sdvnpwao9f2it7NZuqXF/ZU8Llh0x/cQ0fjkCdnncd
nc5XnT912U6IqLcJhXtftYhIj2BXES99Uw56BG5wsWXJnqCbR1fqQJLJUY6MNZtChmCKV84Q44sw
WaMYLMAKHIzMljOkxKec6RQyT+OfOupjxKGqnKVXuzUr0S/Vemfd7+dyC54ieaz7K7SyjjdoFYKW
d50B86ScauQHmEYEpV6fgyIGR/TP9aDQWxnEO+2dKtmJ9N4OgL1VDz2iSF80HYkNG6sHWlrsow1j
Uz/rVT7TSGpdM9XjGRZBVPRDDXLsMS55qBlvLnzWxsMoJoJoujXBhFJe0IPAnXTwGa4gNeFONvxF
yZrRbIDpd8FUAve7xomDYnUFJkWyTuMZI8SSjSJKB1WLJCeEhgRInrmhDhAZrh6YPiQ+g6IeVnYB
S4Voeg+xJUlAITfQmgu06vQWdfmIuM5N4fBnBmxr5VDn2H6AGFHPZlz+Hz6O4WhjJulMrNnhmnpd
mGNzYT/A7+2CiiehpTNSYYG++NFdTAR39ruhUj0mmkjuktCLAnyaciGO35FAaB4RguO5jQpmOuau
RNR2n231BBHLWnXnXSvzlmN7Q6A3dV+w3NeurDSBxzZ0KN77eed9TVRrltsLnt0vyaW4SrZAlpMv
cqmW7YeKOdMDLEQxN1JVtZWX0EJ06WHBOdPUnjfSpHkGX3hseTuRy0Cg+htAFw2mjXlOlPxNQbsz
dienNb1aRvhzQvJH56q0fDSo6Jk=
`protect end_protected
