��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��,�y�}�ǰ�=4d�H���`I"��W�`r���T:tB�T4D�m�)�	1��I�t��
��8(�8t>s)ו�."[�漆���]�~�]��;�O(1#5�-� 偙O��QZ��~rL'�x[�i,mׇp���O�I43��4d�,�H�����SN��d���3���r��m���̨T�I;uj2Y� Er�*p�Q$Gm���p�V�`�2^���,hz�<p��l�Bxt�5��s��\yq���#�@W���f:m��T�	,*�񞭋����_��㧋l�	�\�:��uGd��PǷ��N�I��_����Tuv� ���us�(H�~�{2H�:Zor�Q	#%�3ˠ!��iS��95�,?�.���/�F�i{#���Tp5����Ҥ0{%���2vpn���X�����@l����3dc�ק�3	�Ed&3�ZN O���z��s�yxӡt��v*}ԫy nj#��lc��m戭k[��5)�A#�����8�!�]�Z�s�M���t��w�!��'ÒE�rv��Ϝ�c@<U��\tq+��&|�&X1)C�����r�A~��B�&�����s�:n{p��͠R�X⺂L^��R����c���f��J^?��ܣR�O 1�rV���:��T�4���AD����˩�F�w��)Dm�O�b,�a���1$��c��7t[i2>�ޔ0,S���󧇳Ϟ�ᒨ�-��}�!6��Jyv�醊�^_�(�H�(y^����o#����X��3-�k\8�M�T�"`R�DF6ȕ� �,5�;Ҭ C�k���1\������k�t־9�}���� ���QHF��"��t�9 ?��{E_�7��!����](�S��0�q��w�9��=�i]�1�GʦȪc�W�XC�|�$��}q�6����zf(����լml�dz������*�eLD�*�,�m�]ہ6����D�Gw� �g��' A���FX��\өܹ&�6�h�Ð�$�(+��埧��= Eza ��찠pr[�c&��nP��x�2�TK�M�V���3Y4vIR\������ɭ�1՟?4�_y�y+����ƄJMm����@����m�����c�t�����:ud�Q�����T4���QxBŎ��\o���t�*Z�$�*7<�t~eP/`lfhg��6��[nn��#<����n�D:� ����4�����%=� �@��җ��pԦ������̐z���Xb�L��.�VS�/-�&�~L��c	]s�γ���DJ�����f4���S�쒎l4h�!��>�K��Ӷ��_�+ҔX��c�u����,3��C�l���:k�I��q-��Wb��l
Lr�$۫�'N�0sXA�&�	�[I�iMK�7��7�i��gl��_���� �髖�Y�%mJb�Lna���Ձ�Rb�'�����D�J~P��v�M/���JI�d������Hh�� ����(���m�� ė8Q�=L6���v�W*��H�N}�v��gu����`L����F��1%|���wf�#�0����Q��YAǱ�]6<tYt�8e��l���q�{���#���j�t�_��N�������\r>2�&BZk��P���u�����=.��Ƀ��� �_����C����-�LUg�����k�D8��o����+H[3I�_$O�͜�Tc֘�?g�u7��5j1�P 0�<77P��:��5�[X�U),!�X�9_�Q2��Ī�ӣ'�)=��s �88F��fK�rrK$tmHXw��V�xQ���BSkJBW�T
���L���p9�0����3-��M�I|�����3��&�k�k�-R���٠� ��7jg�R�Lu�!�<�d���I��Yc�Q�<O�V|O�ja�:�d����٦	�����7ͅ��IW�-)O�Xq���L�h�џ�N2�Ij�z۬{��k�@�����p�y`q��1*�Q��Qn���@��Z�B���N�|��~-̖�$a�Íӫ���!u����[�'�y�O^۫�, �_h���>Jjb��JUs_�g�n܎�x�c�Uq^xI[~������Z�g��F>�n|Yj��U6 �r-aR=���@����b/~��o�A"z����?�&��ɮD%0�V�����e5��2[�m�C.Ul�p~6Fd?@f�A��2�/x�^lo�)+�T����R��}^`�B/�z5z�䧛V8�T�6�0������s��Z㩃y�l֙I��I���	n9?�Ϧ�(B�T\�6!�w+43#��9�j��]�[�EIt7��<Vc��jWy�O��