��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����N~@#�k�0!����+��=L���0�ԴZ�2�Mc���ZO�����=�����վ�	"cqw��a��TS[��{=:�����K��-�մ�(��k��N�-� 偙O��QZ��~rL'�x[�i,mׇp���O�I43��4d�,�H�����SN��d���3���r��m���̨T�I;uj2Y� Er�*p�Q$Gm���p�V�`�2^���,hz�<p��l�Bxt�5��s��\yq���#�@W���f:m��T�	,*�񞭋����_��㧋l�	�\�:��uGd��PǷ��N�I��_����Tuv� ���us�(H�~�{2H�:Zor�Q	#%�3ˠ!��iS��95�,?�.���/�F�i{#���Tp5����Ҥ0{%���2vpn���X�����@l����3dc�ק�3	�Ed&3�ZN O���z��s�yxӡt��v*}ԫy nj#��lc��m戭k[��5)�A#�����8�!�]�Z�s�M���t��w�!��'ÒE�rv��Ϝ�c@<U��\tq+��&|�&X1)C�����r�A~��B�&�����s�:n{p��͠R�X⺂L^��R����c���f��J^?��ܣR�O 1�rV���:��T�4���AD����˩�F�w��)Dm�O�b,�a���1$��c��7t[i2>�ޔ0,S���󧇳Ϟ�ᒨ�-��}�!6��Jyv�醊�^_�(�H�(y^����o#����X��3-�k\8�M�T�"`R�DF6ȕ� �,5�;Ҭ C�k���1\������k�t־9�}���� ���QHF��"��t�9 ?��{E_�7��!����](�S��0�q��w�9��=�i]�1�GʦȪc�W�XC�|�$��}q�6����zf(����լml�dz������*�eLD�*�,�m�]ہ6����D�Gw� �g��' A��)�m���b�����L~�B�3A�/15�s�dm�\��rbY�6�g��x��E����Uf��)
^fd���YaŌqa���h��!�u�V{�hPKS�1�J����>+	CK�Sb�} hS���y%�Uyf�MW���BE��=,"�L���Ǎ5�s0A5��E�)s��O7^�]�Y�٭2�,<�>�]`�k�b=!�!����0y�k����WU�}��0��(-��I-ip ��J?�ċ����j+Q��zR}���K���a�'2}+�Qp⺅��l�V�`<AxH_��P������")����7��cR�8�����1�Ϭ,0Ê�J�ߡ��� �B�7�4�q��#Ddۖ*J�%Kи�ޣ|6���hE�K���=n���"��Bߔ���[kAT�b����P.���c��5��jL>�m%��B���n��y�r+�v��+^$��ۅ���U�ǉ��c���3Kp�l�/�+=.�ߩ=�D�"�?o8|ޔ�vv>FЫ�
0j��B�a���=��8no�a �J���*�#?!��4�0����i ��'T�	��H�I� �EB��,��]!ȯ&��,A�O�F=���K���]�oAy5�t��d�O���s�]����X��g���;��r��hO٭�d��\���l�P|V��u#"+��7�H��=�?t�Y�X4�~e��1���l�Шy&]R�F���BNĞ3H����*:2_����7���h�2l&�A���%�l%�Z����D�y����q��"�Mq}ay�(\!�\௚rj@WsX�Z^�m�7F��`���ae�9�<Ұ-f�D��*�D��3d�<6)���O��۬]jB�j�9b��ofe��	5�ڣ��,$�u��=4=܍ʕ��"�y������]���衢I��Q>�#�ηa`B?�F�w�ɿ��L`��>�C\�h�M���Z(�'��M5 j*}ȟa5Ͼ�PJ�W�WgwA�>�c�N��i�$����p7<V�b2k����_�r�@o��DSk�:��h���<_��Y:�k��U{=�db��2��~g���({�&Xu��ҘU��xtwm���=�{,[�Ϲ�H�_Z�����
�y}p��r�Ȃ�w�a,F��)N���a��5=z�:�P�����r��v���V�ï�V+ʟ"��	�#;.����:	�\�Ė����2�T�cwЗ�6�\�pH5P�h��%:��P����=��b݈�{���&��\s�d̍�B�s@��Yq�����r'Ov_Η��TaCf_2��?E�+������cHS��~�nR�䒁���i|cX?�~(��G�ТRb���O�<NN��yt,z������a�Ѯ������.�����KS�ڂ�K�xH�����,�ݭ��(خ��5x�is:f0��[�,�>��6i0<��=q�x��:�e�%��;ϡw��d[�1_u+y)5n��)s�ҭg"��
���G��kR���1�r�����a?q!z�Y2�:Rڼq*�}ߟ�0���+��s�?�����ն=�P�C!N�&W������d���ԥ��La�wk��|��%I��f��"O¸�AQ� W�-�!�h�I�1c��}��姙t�KYP���h���1��zm7'�[���N�ѵ���Kǒh�t�7sx����q3�BOKG�٦w:k���@hKZ�6μ��|�M/ռ���8��,�c�|"������2���<��X�RBNu�e�-�^�Յ�Q_J����`1��3ͅ�+�O�h6�1�U��k�/�gUmE�>�s���V0����NT.���E)�����ð)����k���(l�W�� �G����s)t��I�Ns�O�Ga�>u��	벒���y�����W��
���'ț�Wa���O�,�]j
� .`�\�}s�r�������o%���H����
���j�T_�U�.h(>]�2��#w��!K�-�7�R�ޔR��9��F�)���Zc�_����F�āTp�c�_߾�z���ö�\��l{{z��4Xڽ=:��P�`f��	�W�Z��-6���8���>֨�ն��#a��~K3���|40�������w���o0��#�� �Aj���f��3dv����3�y%�Dq?�MN�3#<;��^��Y���(�_\V�Ϝ�)�[�f(�i��C
Q�2Ԣ���>�>����}%��9(�B��|A��I4�5�����*�9�zf� �p9'�^�ƪ<Z�Hw�$� fL�-=�i�mU�q6���6�2O��9!s��%��𝘋���B����#�=���{�U�f,�4ς��.��<,��_.��^MgA�(c��p^}�S`ez��e�j�i��uX�����/FbՇP:�(���[CY���wA���+�&
ψ��a�4�m��A?T7�� w!F>��-`��kgS)������Я�X�� !S��U#˒�G�=�Y�}5M���2���H��&б�h�@��Os鈣�r6��~y�,�r�@2
;b�<�C�Y��إ~T��d���-ĉi�%H�1*?�^�V\_ ԅg�Dt�"���$Ŵ%,�G.WPt��X́���˓[|�΃݉6�~b$��)ͷK�|n�.����q�H�+��8Y� C�/$��翡@;���W,�̖�TZ�z�F�d�~P���ߺbT}9���gG�o}�F�cE����崎��+'Q�4�74 v�F@��&�KӰ������)�Ls��� ���㉟��)���˵3��l���V�����p�Dġ�qj���eu'3��[(y@f�S��WD|@���2[e����sߚ�*��v�l���ɷ�M�I��s~������,�	�Ҷ�o��]����P�Et-�J�o���c�:�"āS�Ww����>ѧ���@4.8(^E�ι���s��ӋA����g�q9��7��h��]�ϩ�tF,�U�M[J2&dS�+�/�%��dD;�xk�A��.�xx�*�f�<WL-O�j����(gќ�8*z�P�ֵu�������C�lW�ɉ��T��P��@f0��X�O.��L�����Cq�Xs�z�7�Cd���w^�N�U�4Q��S���*�.�L�%�3�\Ƣ1q�|Y9��	����ݔ;Ȧ�>�]0�Ѧ��m�.��o߯iQ����՛!:�k���N���9YL�1"O����D��0uR	�kk������4XJ5_�?���Fl��������$Wj{�k�3c�w,�읠�%!x<s��3�|��ˮwε���J�.��5��A)֥��Q�9衵����"3)��Y�~j]�fR�
֓s1�A|#Ĩ�T8�{�8�4nVrq�F�QW�F嶾�={a�ߞ��<w0�=��&bɇS+X��Ų��L޷l������feR�6�>5Z�hz8�mW,��!�\�ơSy���)6�N����s���XJ@�نdcf}��4�6P��W�ק=�äL;��ۆ-g�=�i�8ri<��`�E��|Jh���e��0�-h�Q0n,]� �������N	t����޳_B�\�_k�О�������d0�y�Z�i���Q��I"�=uqUlXg�yJluh Ye�Ś�a_���"���hZEt�Vۥ��Kd.r��w���Fn��q�
u�� ]�e˚���:�+�G,�Du��*t��2��a��*����Mv
i�G��y�����m��Ϩa��dý�b���C��*~����^�/`U~��d�!{��_`�	�;3.?��1���O�7�t�;��a�9�E�����Q��w��hR����?��@���\�[�$��)�Þ�}5=s�f�����J�s(�x�	.�W�L�����R��(q>Q�D��6��F���f�b`hV�U��L��<����8�h�J<^��Y��i{+i��c{'VMk
����I�G ��Bλ=݃�+#m>.�%���cIN`u�(���
aL\HU���-�X[�?���nO���ym����D^�:V�9�_�>E�]�<¾%{��e�u�Z{�d5����Ñ%x����Jx%�[x��e�5gz��7�z�! �x˃T�K���'�����B�Dq[F����F��V�D��$�\�2�zU�+���e����lB�F�D˄��#�G���Y���F���1��H u�D涱��3�=~�*0�J�}�&��s����qЖ:x�����p�<�J��ś͖pPM�S9�=־����w�l/?Ƒ$x1T*��n�h�Tf~Ɗ>��xs���ɿ��n��ݚX���Z%�h|-B �<x�0é��F>�G�\������G��M ��ʒJ�A]�$ɋ"ǰ�z�?���{:Z�P�ͪ���T�u���Rx2%�}ݻ��_�ǁj?�ԁ�X���En�������{����sQ�ᶬ�� �
�S�gU��j(,灬=���b��FI��N��G���o�~��3&����1���6�_���ꙫX�{'�G�T�m!<���2�U1yo��5��R�'}�I5��g�%����7 �{��������3g����E{t�Ѻ�TZ�^�2+���]��:�-�Z�!�ⳁ�c�|r���Z�� �<6���fQO,�~�^��3dݞ��,���j�wz�=|��0K�����KF�`�,2J�Q�9h ��2KԱ���,4�n/ �ݡ�y��G��KP��G�#�9MG�|�5������Y��`zՋ�r�Tü����7m�	huZ������m��	���3:�K��h�x�(O��e,\�ҚO����ė�����@��!7�(7�X��-�[ʌ��r�# �*��ьDJ�<H�ă7Sg#az��k"�j�Yw��h2-��%���Y2�����gWTj����+%��m�.�(� u ��ˉ(	��>hn���4XQO�����>]0IFe3_ o,�6'����3��� H=�O"�
�(+���Q�9��8/_Ԑ��/Uέ�'9��*q��P�</~�8�V��׹��H�9u��]��h{n��A=���K�M��)�Pg��	O1�Y�/�
B��W��z��	����ꨱ"�o����%��_F����'"�ȁQ�\d�3W��t�U��6��R����A�����ח���_�t�E�
��o�;�u�8B����4�qOSqDO
&���QA����EG~F�]�F��aqy�J�������먑|,,v/����E��s�͖��i%�S	����T���4��F�K��(S
"Y�F[ܸ�|q�G��z�ދ�8� 
�4���_C�;�V�@��"uy$|�-�1C%)����ޱ�z����ܳ�)u������M̫
��Ȟ�s8�:������{a}�3CU��>x��������m�W�] b���1���[󏽢ƺ57Y�"6S�j��I�N�`�̇��h�W�Ƶ�:���1����/d��Ӷ)�����)[&��k6��T��b���q�n�/'pz1Y���ƪ��:bRf�n��ՙ�]$
Ur�?x}��~��a�
��q�{/�M��|'�g6x� =m�,�X7Pn�:;	�I����}���b�nE��(��Hy],� x:	O�m���ﻷ�ˎC_nd+=��k��\m��n���[�?�`��@�9^R�x���a�Q㠧#��k=���X0q�"]<M�.�\�&������*)�{�0�]�\��Lׇ���{���t������c:��\��W��1�
	\QL���Z��D�}J��yP[ѡ����"���@_��s�fyPJ�]�׈[����M�F���>��$ �	4��"��X`-��~���|B^l��C�,�����7�+���g�[#��D��y-k|��	X@�V��)Ջ���48Q��>�`�#������c�"�;\�zEЗ$2r����`^��+���q<�����y����)~�ջ�6G�=�0��ì���r�.۸���h��]Q�����/S�fg=N��VM!ƚ��,�����p��B+[�^�~l��_�q�s��8,h�����B��˼��y8L4��|�+��CC	��1S��35�^��L����ٳ�h��| ���J��V��n��-Z��&Cr*�F�����N�C�)��Ec��B�Jc��_��(AJ&0��̮A���x��h��c�)oQ�p �����)��Qt��~?������sn�D̆�$}zp�\�̬$�H#r3����n������=�۠;�{+�3��Œ)���P�5�A�$q�������-��b����Z�#Ϲ�j��o<��DN?����c�Lc<�l���Β��1G:������ 53˚s՛��y��'���^�<o���UZP��a�  S��&hL�<(ECo
q>D�FH6�߃<�@�Z) R\�1d@D���@H�(݇����-�`u�b���o�=\��\/�b�[Q��1|z;rsۄ��X�6\GYr�{w;��-�S��%��k�>�G)4��R�'�� ~L��צ�3;g����#A�R`���[0��/�B&��T�ױ�����}2��ѭL����	������I{m�����c����7�aN!��\�7.ƭ��L�#}䜳A��~?.�����~��0�[�p�@gp�3Oaa���1��H��F62�l�������0�U-?�#OFy�*�L�]�w�Ž�l�&(��\���gY>�E�����'��aj́��J����ɬ�u�$��f�P�0�dБ5d� �qP;�����c��gW_�
K-;�H��8��I T1\U�^S\2]���'�Wk$ _��|4�E�m��5�QS�֣`�ibk�1z�(U��V>0f����<���<��G��>����3��x.B`��ɱ$'uȲ�%/T��4q��8VD,�c���%'[�����(i�q ��:��X���E�}r���AW�t�K��h�
6��O;���i; K�f�ώS1�����",�<al�W�/���IqƊ=�!�.���h�N���&c䳚��SP��f���b�'���`�+���A�)u.ؓ^�4�Sh�Ug���4����Ff���' �t��t~*0*����Q~p�TX�h`6E�p|�����Q> ��x;d:.FU�X�3m$��E�_ņ��Z�7��m<�~m��Ա��"�aĪ���J���4`ab�������w 6���，�to�5%j�SŅ�D{Pt���إn?�ȓ,���C=X�Z���.p�I�G!|�1`�W6(Kw��"�Z��
%�-���DhEoՂ[�#�m�g��P�;�U;X�T~��d`[��sX��ߕn��%�;,^K��9Î��Ŋ��f�H�̓�Gp��'�9�7.����I&t�<�(��e��#PxW����(f�f)���1�v]֍5�k��w��w�-�raH�#��Jw~i@�p�'�(ڑ����k�����[�r�)�ʼD#^��4�$;�(���>���7�-�P��Z4�6�}F�K\k�����d�	@R�,,� ��3�T�ۘ$����ϣvǨ��I4Q��U�^6e�f�Q��n �K��PQI��{�}ޕG.6i5�w��8=)�8ⱹ��	q��9�5��������LJ�̐;em��U �$���4x!L*`Gq#