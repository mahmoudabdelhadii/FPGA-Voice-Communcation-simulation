��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��,�y�}�ǰ�=4d�H���`I"��W�`r���T:tB�T4D�m�)�	1��I�t��
��8(�8t>s)ו�."[�漆���]�~�]��;�O(1#5�-� 偙O��QZ��~rL'�x[�i,mׇp���O�I43��4d�,�H�����SN��d���3���r��m���̨T�I;uj2Y� Er�*p�Q$Gm���p�V�`�2^���,hz�<p��l�Bxt�5��s��\yq���#�@W���f:m��T�	,*�񞭋����_��㧋l�	�\�:��uGd��PǷ��N�I��_����Tuv� ���us�(H�~�{2H�:Zor�Q	#%�3ˠ!��iS��95�,?�.���/�F�i{#���Tp5����Ҥ0{%���2vpn���X�����@l����3dc�ק�3	�Ed&3�ZN O���z��s�yxӡt��v*}ԫy nj#��lc��m戭k[��5)�A#�����8�!�]�Z�s�M���t��w�!��'ÒE�rv��Ϝ�c@<U��\tq+��&|�&X1)C�����r�A~��B�&�����s�:n{p��͠R�X⺂L^��R����c���f��J^?��ܣR�O 1�rV���:��T�4���AD����˩�F�w��)Dm�O�b,�a���1$��c��7t[i2>�ޔ0,S���󧇳Ϟ�ᒨ�-��}�!6��Jyv�醊�^_�(�H�(y^����o#����X��3-�k\8�M�T�"`R�DF6ȕ� �,5�;Ҭ C�k���1\������k�t־9�}���� ���QHF��"��t�9 ?��{E_�7��!����](�S��0�q��w�9��=�i]�1�GʦȪc�W�XC�|�$��}q�6����zf(����լml�dz������*�eLD�*�,�m�]ہ6����D�Gw� �g��' A��)�m���b��ӎ���o�6ūvO��=�W�������}��	����z
��z�&�P�K���Fn�kU,{��:Ծc��%(h�=u�ݦ%��t�|+ǆB�������0�yȒG�좩�����h�g��M�����!v�+���#,F��iS�5~i�� �ؒ`.�|NT0h>�~���M/%{�mh[����<ljd���P�Тi����F�Ϋ���g��j̆g^�k��k����A�s�ہ?�%�C��;xd�ǘ���.!A=K�,K�9�>�4�4��[�A����?6��gS�mv!����0͘��!��-�,��Wr�>B�|��n]��c���]�r�������ӕ�1�
�;����ߛ�b�%�\��#xg�����zkד/�s�>K~��������j�TZ�u����ۢ�PʥWHK59Օ�,�]]�wg|>o߰q��
��#zg�˛3�T��x��2Se�K�i�J�o*	n���>�h��e��pβ��� �zZ�8����9�4}�s��ͦ�D��4�Z� [������lѢ=���&�����Bl0�jZ#�����(�=����b�lL�@�^����)�t��[�z���U�p�9��\�ºH,�!U�����5
nD�Nߴ4�u��𡬬���L�u;{���9 H���T]���yI6I�;��G�d�\0:0�q˄U����k�W:O�z1��
 P*`��_�4R�0%ZG��Tʐ��Xkk�����"�dԣOS��Y�J�aN�#4-��q� ��"�?B�y�	�T���9���c$�(�v�?S5�e��1^[�e��u��b�����ޞ�G}7]��SI6�ݏ����oQ6r�m]8���r�_~���0�^��:�(���nr��}�A�{^�2�.����_��֗�X��2`u<�ԉ����u���[4���2[o��V�)�y��P=���\1�O k�`������.0�&��?�e�\�e���1�ܹ#��K����2j,Oj��N|Q��ic����H�Jp��LJx�9�0@�%�Ѡݾ�{(
.z�����*�hH��SA��>�Cw�w���#�Q}S����"��/P���L[��������Iv�^#eN'��|�l q;���(�;���FZ}IW�+z=�4, z�,�xD����vD��/�F��ރ$�s��P�=G����נ���V���v ɏqѼ��`�*�׮����LD]�6�y�쒦@؏7����Zާ�2��U
Z/��r|ى���%(V���S�g�|f�{��s��_r����W�x̧8S�&�YZCG�����}�ث2�YP���1���d;���Ō��]�H��~�8%���a������'��	�fU��؅1d�P;�}�i(�٘ҹ O�� ,��8�BV�g�jh/����!�H%;��8��v���1c �:?_��M\��-=A>�ڙm
ª��u\��*�A�L�$5�P��xQ�R�y�v�'A~P<����*�^�:<&�4���Q|�����m[	\��e$�;Q�~ 2�֜���<����$�r����6Y*�*�&�k�{�rL&!�N���򺌤!�4�r��|���t�|�Dƹ�W�����<��YC)L2�@�����v�S�ţ�U�5w�U<N�D;�^�X1���� ��D��y܎a	h;S~�k8<��v31��w�ԕ�]<�.�~�o���]�~0#�1���ǆ`J���g�g[�^���M7����F�Y���ж�P!˛��\����50-��{��[�0�A�c[�S��Ĩ�}��0pz��-
Qʞw*(�V�G�X��_o��������}���<�6&u4�u	-k��@U�+ړ�ɨ7�����Y��NU~�S�+���!]"��I?֭�H��Df�ęz�ro�g�Vq�Q�l0����.�툫��W�o�<��C3��#z�̇�h���[����G�f�e�5��?S�O`�S�By<�fN�?C;��ʏ@n��ǉ�?��'PҶ�J �!�~��W帷�K	>f�#��"��HplZM�R뾆����6���\�m����h�&�#��iV��P���,� ��V�� 鄘����v�
� PVQ{�_� ��E�b��r�m�7ܦ@\J��+;*&B��r'�@�3r[�	��h�$�����*����� %���8Qf�v��J��<���.�r3��z�zʹ}\�}��VŲ�L[[u��
B!�W`d%�G[ݯ��`�<�0�]9@�)��	��C�Rqn��@�	h�$�,���b�$F-n���:�k����\j�REnʐ��+�B��yf�隣# b����
R����N�yD�y
5-#�������h�B���1N�-�3#�i�r���)"�9^�c8�-����d��F�v�@̳\Y�{�2u;s�a\J�rl��N!���;��<�R4m�.y�G*:�4v�F�A�K�~��_\�� `�X�|��4O}�c���H-d��Hkrq��U��������(pah�̈0ޣ]ϪXi��
�y�E5�k�e��קɥMj�5t�o�@�����>�x4ڇ���-�k��U��������Ssh��E����-d�����ʒYĝ����ܟ� O�v�����&�[|3���ዴ�����K��(�����?��>!�_�������W�f[�L�ܑ}��{;�����=�����HT6�ݞ� �5���lCo_t�'�r��K��Cp�D6h]���x�.�zŕ����,�p�|��u��4`kg�!�:]����`.r@ 4(�������(�͞8���(���V%�\u��arʭ�jG�6��q(������I,{�s��#M�xsW�M���F��''���o�3c�G\�����P���VS:>Ԁs��ҁ;��!�k ����S:]|La��%A	���V�5�p�ɉs,Aid��7���,�Zʸ�VI�5�UCp��[�PP��J"LsM �b��׃7&������Q���L��#I}�j|��Uj���J�<sPq�.*s����H��ބ�C|�������y,p�ի!!X��+��>��ŕ�y��w659��і�F�;�3��#�����l�����՞����Q����3#}.h%���H{�F�m	�(:�mN���:4ő�v�}d����kY��%��3�h�+����#���E$N�&|.�?`Rs��Ԉ���Pˌ<Ǫ��T�c�rE���Q�I�s03�w`��h��T��}��Լ�続e2O�N/3��Z�^��z��-W�U#a����1Y;�P��^@�/�Y��z���N���c�03��R���~���_�� =��n��U��CDl1�Y5�U�c���4o�����;���պ��<�� �6����
�Te��6�f�F*��c�����q�-������Mү��A��j��j �,�	B��s0	�s><RT�� B&��y�'J9���]�kbL����J�\���s��H�L����35�b��M�3k�  �7<�=ގ�T�Gs�Du�F~^kO��Q(z�E�$-KG{�����tWV��;�I eh(2�5!�7�B8���C�Y��j�SΨ�sP�ֲ|�Xт��D�z�a���%���ډ��:}��V��("�_�'}��Ws���J�R��R�)��4(uQ���P��ZٟU�6�gL��5���ħ�"��5R�te
�.����E��P�� ��Qd�1@ֈ�Ѥ\I-t(�ނ��
�y ��Ł��HPV�<_��J��#�<cK��G)w��������+Q�+�!�&0:MH��S�XXN�h"�K�U ����#g�%��4�m���Y���Ð�`�q�q?܉<,�m�jTlkz�������x��f�@kC��]�ݰ�{%9R��I?�ǚ@���.dܠ�	/�����G�Vr��������0Λ�D8�Cg��vġq=�����������k�x9:�EV������7�9]���NM܁�3�3/+!�*���&:��9Q��Z�oۑ��ˀ\V8��SD'>a�#)��x�+z�OS����& �������#m�IH�C��]H_54i)E6zD���꘷/F�4��p���?|	��úC��O���s��vCd�=P��$���Ϲò�g�3���њ_>��4������Fx��'1O� o�{���x�{*���*x�����H�NJQ�� ����C0]qd�*Oa>�/up��䛏X�d��l��݆$e�e�&;W|9�ReL7�̑��;�N@�j����[��]�{`�����f��n�z�k���,.e��bn�1PVK�]1��f���0���L�Y �����j'�U#��������Ihm�,7�K�E��WR?��r��'���a/�����T	��>ڥ�"�)���?^d��7�\;~���m�ð!��z����m���4cS��������,���@ϖ���yj�چ����%J��$��/O'��;O��f����J
��9>6���m6p��#�����$�5��?�|��V���AuS/A�@[c�x5���݆��`�N��8��%ۨ񃄢��E��w��)=�*7���t���mb��D+��C�2IV}�$!5c59C*a���S?m$�@�sA�����*���MGW�LA�Y�zI��hw�=�\�+�8;�B����O|�!� 52$S��k?,˲6�W��
�����8�����ӇąkE��T5,=c@YOk�V.oy���+_��ѻ��J�rq*D�a�������UF�]�ٙ����7Y���4�u�q���Z�v������5�l����D	��=����l;�嫬����-�g���6��}�N��K:9�ގQIk������X��3޳+;[F�MP��c�X+ ���%�V������*:�9c�C�*QDM��ٻ�{^.��ѪQ<��^��/%�r�����D[�G��]��Z������9�}�E;�?��&������_�Fƈ��f5�=�$z���ު�j����$�[H<��ShF��*Nhcl:*��#a��3�v�8q
�GW�0��/�c]o'7>�v����-�sE�w�i����6���}����C�%F�H'Z&��j�ߥ0��K��R8��ޮu�rꧤN���# �HD�iV<֮�p9)�hyȔ0ї�*���_em5�L�#��nЊ�\�ԌO���=�8 x��%9S��D�j��
�3�1GZA#���>a��Z����]��p�n��^&;��e0Q ����|yH'�"g����"3�E�!�[^��Sv�)��n��P�J�����{Sb��%��� ��{8	��ļv�:E#�jr��dY�V$p�Jz{�kKј���_�t�J^6�	�b�n� �o\A���~fB6;ED��<x�R���ڜ�8)���N�#�t�4?T&doz�� ���'B�U��@C̦�-�BZq��1G|�%/
5!e`��fLFdH����qJQˠۮ��/ �,^IxVSdiE��d�rU~�UQ���0I-rS�kga�m+bԞ��M岯�T���	��N�G�{�lE,�ɱ�������I��w���r�%f�|�(@[�W��%�E�2�Q�.R-�M�����<$:����@�;�ĽWTk_��7+4�3BA�-1nk���oej�pD��n02�kyA�L<�NH�ڄv-@I��dxT�M��貨,�4,�I���"+�[6?�6�f_t�+�$qbmu%I�e� ���$��T<@V�r�D}ݱ�r�"�B��$�c�Jr������{1so�� �V��2�ߛ~���:.�%�
Qn��'B�3�����Mw��2w�3-U�ڽwr<��#"���J~V���o�R#�=�oY��=d�����kWC����B��HNH�1�a%��]���f:ێ�z������1��1�~1�T��
�j�e}_�[�>+Ǚ�X��酒:`��Q���3�)/T�VոL��R�Fk'��qOF�e��w�R�R�S���>7���j�^no��h���N�~��q>���el�vu�u0�kvq'A��9�{�3�fv��!���8B6!����|�$+�_Ъ��Y�xށ���4M�g��@-�1
�J���"�}@y�H��a���!!3P��[-�{%�$2F�Ѡ���#W.��g��2oji����Beڔi�Ap��f?O�(4Qf��-��-*�a,��p��i�j��n�]�q���C�.�t���-c�/�[�ϴ�`��$��Z�~jT��Q<�qz0x+5����
�%6��� :�Z�����_�,���J\��U k�s��i�$I1�0�h#%��8����A[��!�|��z�k^�x^l�A�|��Tu2��y���%0������c���I<������ar��A��@(���Ǿ�^y�,^��h&�����¾~�4u�Q�	ښ�����kơ*��k�q��pa��đ�Ā��b�Y��̡�3�M�ɢM�>�2��i�L�g:�^$h�*��$��M�yB5g�h�])��V[��k�p��"���� |-u���W)K��%��x?���a k?��y-�.��i�L�������6�{F+>%)~dC�7���o�c���?I�|�ʱ+�&g���\�8dN�}𿟞��4.�X�HH�o$hg<�^ X���c�RPNH~�Q�V􌠷�
����Q�"��d����־/R]����o
I�z�ߦeD �����%���3�;���(U��a-���:��q������bҕ�~ۤ9�{�E7ӑE�p?�KA��#~4�,�k�d�B9h�c�F���4nV�u`F�+�\�s�3�/Z������7s��xa�z���?��nu#ӕ���1�u<s*��D�y��bC��p���!%���,UI�+���C3,l����;�+.�Y��Y'O0 ���v�s����8�}�!dۖNǁS��7e\�7Ҭ��+��\���^��9:p9�k��˼���]�%֠�����arz]v����厴��--�^Rt�t #����}K�n~-e�8>��
�h���Q�v�B��D�S���Jj�@XH)_�(C�WEW~;��O��7��L�����W��vp�``���C�hl;SN2�~�xT��Ԃ�DNU��uN��ɀQý�����ɅJ�+]� �μ�}��k��|�2�{�}c��քk�Z����.����h��c��s�� ��UO��oHl�SU����O���(�����9���S�����y��[1L���^�?��!�u�'�������0a#�p:Ö	�q�<��W�Q�x'1g�����D��l/k</��V��:��n~��?6�^t��g�ׂx�hs��`�au��շ5��J�x=��,�GL���TJLΉk1�ۭ!�h�M�+e�	3,~��pj�P%Yxd�=��oJ\Td��%� �joͯE��<��cs��� f�bLW�6'7�Eq���4HM���/>�i�윿 ��O�=�����p�D��܈���!����m�'z�l	�o�'��c���8�G�c��〿�;7zr�?#`1�����wt|��AvǳgrM�SjR��n��ze1��ΞY�-`������z`;��,y�)[xo�6�RK�}|�������<��B����yQ�2}��-z+��Xfy9q������uf�x��b����<o������!A�.��t�}F�U���s�gB'C���U��*T������t=��_��j4����K�+����î�������Z�+~*<(* YQ��WX�ٵ�Y5����n���K4_�P	~�W�!{yb���rC���vP�7y�9�$����r�������坻�/�JB{d�	������@���
�h�f�GD�+�q>�&��į�	?7��!�M�Q��BMO_���e$^�H�;�)�x(��x\�`em����}����M��f������k8� s�0��v�P��:P�=�nU�x(Y-{d#��Y�4��d���doVOt�CK�a���e*aT�
J���*���$�*apA���o�J�E�XD
S;1^4�#��e�U5�q��,徰��6>����p�`��&�,�P����N��m������5j��S8[��gdO�Rka�P����5�ni����QfQ
u�M��C�B��H��U!@���s�dp�����G��\��OW#�[,2@�@~6p����&'?� �k��&'2�5��<ي��B������d���r�5Pl�0�̗W��7��Q}
ϸ��MF=|'|G�\9�"|*4��C�[�H�P�'�x�� sA�n؛{�-0X�X\g���lG�U?�����,6�o��v�/�@�_y7�~��tƨ��;����i36�%����p-f����7���f��1)%
j���C��� ��p�c_�SExr"04��q~ ��������F��1�B���3kA"�l��S�n�ݲիm�J$`�o�vNZ��ZP�n��ƥ�4�%�	�^�\�"o�B�y�t!�Ή%�E�׎«�΂�)	C������7��1�.,Rߙ���MC��lz�*I��1�sxe� 	���I�D��Թ���'wL5�|���KӪ�#�ع��K�8�z�������X�3񣬐�;��0�s�Â�bzc�"yv��>������s�ZH{�����\0�	%���(���O�bdԞ{����b|�A�.��v!zS"^O�Kn<��w����8�� ﷴt�	LU�v6�O�eu�T�YSk�����������x ���^�Ռf���ۣ��|�����c����я���Wx�Ey{Ntp���hŘd	��<>kb��������@`���'��IW[�!6�xu:e���Д,�S4f��ͬ�%:�_MU"�%�Qi`iY7�"�z�X,(VN,�	�ZF���5�RE���S��
����	���~�̘��_h!����q��lJ��mD��^krD��»G���!ɶt ��p�?��c�j�+�o���8^���N_~Z9���y�}q~�5ң���-ۂ��#"�Ɩ_�/��K��-��@�б�3�22Ӳ�1x(��J����|4�GK�f�taC�9|iy��
��B���R��Dc
C�n/��
�3rm�c�!��q�4�D�q��ub�7\ӟ�6���Z�-���n%���m�(��y��0]�?�q�̂�ɷq�=�U��LW���|�ܚWV,�{*�2y ᝱	7?JJ��ܔ�[.6 �u��`�x�}m�5���f[!�H����z͏�Ӵ���K���eз�2z֢P �������?�_�	�6uOΛ��v"2)���oV�:{Iu+�DA *<W����Hvk�ё>ͮ6���L���%�+���-W��q�5��c��x�[��ǙlX� -����8���rL۩p[�� ��UՐ{zt�R�$����{j{=�I�.�u_%O �z�������A��#�
��[_�48�,�/����������F�O?5�UI�p�[I0����"j93�se\u�'�QfO�9�w2�-�|�M�K�f|�U�5 ���<��C/a���t�B� ��8H��'W%���Ko��o@�Wߝt���%�"���-1!�!��a�"w�s����l�t���+ݙA2|��t|��P�P���7���	iY���+Wi�R���q
:���ۺ�-g��F�g�AB	�>_�5��i*��{���-���V�b `a$`l+Va ���s/DA��{<t6@gW$��J��ż�K�Vj��ki}���{F!m>�F�P-��$�J���O_6V���4ޑ4P���X^!�5�]�i�B"h8�L@Z�n�8�K�*̔���@��=b4Vc"X���N��ò�[�w�I��u1��ۉNueR�D'�7Y���)��׵5�����5 ����ޡ�}��A?��PV��n��0�X�q�^��?��u3�'� ���Zs�gE�V
���厘�+�G�Ќ�;��y�e��%��8N�>A�AXRZH0�1�NWU^"��M�(�mV9d��|�}���L�7wj���ӱ�:���@�C��,[�`���pf��,��F����(v�%�uą�����fȚ{���|Q;�t��=���v��a�W,��d��>��E>|f�[gsz�b�=;���C��T��e�v=����[���>���.8@�x3�d�q�2��"�� �`S}��^�p��R��	�v�叉o�a��O����	Th��%����_��kx��_�M��nz�]9�Ҟ10��n��f�;gз������>gZ�i�9b�P�\��X�E��RB�L¨�l�-��z�5�o����)J���j��Q+*P����z�T|l_�ɬ����������W�����2�E��P7wЖ��<�(���&��qe_Q�'v|��-�Ab� :�k�XVtU�"��v$��]J�����\ʳM ��l7���z��s������oA�	���M9����G��2a�쐦^�Ǥ
bj!�~,��S�|�6�i�*^�kz��A�xԊA)��Ԑ��c߀�\��/*�Z����:��֓ɛ�EшP�n'k ��d�vde}���-Ky̭�mP�n
lw~/;��C�Vʗ�[ߑ��MyHΞ�#�]��F��l�xf,DH��A���u��	[�E̉���~��>4�N��l�O�3��i�1Uiiª��ݷ��r�$��s!��`��^��u�Bt�تm����$�b�6��:d@h��r����F?��r���quF�ٸ�.@)j[gU�~��g��؝���4_+����C�,(	ʭ��k~0 ��@Y�g�p��6EH��W�kQ<ݙb��GBb!3<���Wf��"�H��*p-��[S���i7�}"���\?�֮u#����֫GZ��e�.֯NS�%�y�^��St�2�jK�h=Ca�J�p��C�h���vW�@Y�:��WB�i�wp�N����ZE�E=0�?6������j#�ܐDLIS��*��cdJ/� ǚ����T5�:���#��3a�+ȃ
�
D�~%ۧ���BG����L)������);Tɺ{������ �BG��A� ��bB"<��r�XV�
}bw�0�Q����u{$�v�Z17�	6�/1��{,Sr$x�	YY �k\���w�2�ou�!q�x���g�C�9������?uD\�i��5��gOdE\}�U��ƟZM�7_f�ǞqrT���ol:�jp-���s/b}�Sˇ3�L,W��0�Y���ް֛�̚ד���3����b�YR� v������:Qg�4&�r��g�ԧHώ=%ԏ���҃7y�,���t{����C c��WXA`��{�>J�rרSPV4� �V���3��7b2���YP&��z�S`�󚙩MV�#0�EEG�7���1����8��)mg�"���!θ���J�K��@��2����N�0�Ңw6[k�X2i��%
mG��(K��qdЄJe�a$_�$(�Cb~Q���R}��$�u�R��}��vNYL�[�	�k���@!�q�<��%���ʶ<�*�^����d���XNi`'q��B��� �"�
p9���	�p���K�J9E�",���-EF����N�+T�O�P������?��*���	��[Aޑ=���j0���1?�[� ؟��G�C�~4�=�U�Yoh���+ů�@�zDq9���W��`Qx*��o˜WU����z�(��Z�P�aM����xF��I��s�to�k�enK����ǒO0�ؤ���c�;sgy^�Q�������a�V<����������m6�ꑾ*q