��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����N~@#�k�0!����+��=L���0�ԴZ�2�Mc���ZO�����=�����վ�	"cqw��a��TS[��{=:�����K��-�մ�(��k��N�-� 偙O��QZ��~rL'�x[�i,mׇp���O�I43��4d�,�H�����SN��d���3���r��m���̨T�I;uj2Y� Er�*p�Q$Gm���p�V�`�2^���,hz�<p��l�Bxt�5��s��\yq���#�@W���f:m��T�	,*�񞭋����_��㧋l�	�\�:��uGd��PǷ��N�I��_����Tuv� ���us�(H�~�{2H�:Zor�Q	#%�3ˠ!��iS��95�,?�.���/�F�i{#���Tp5����Ҥ0{%���2vpn���X�����@l����3dc�ק�3	�Ed&3�ZN O���z��s�yxӡt��v*}ԫy nj#��lc��m戭k[��5)�A#�����8�!�]�Z�s�M���t��w�!��'ÒE�rv��Ϝ�c@<U��\tq+��&|�&X1)C�����r�A~��B�&�����s�:n{p��͠R�X⺂L^��R����c���f��J^?��ܣR�O 1�rV���:��T�4���AD����˩�F�w��)Dm�O�b,�a���1$��c��7t[i2>�ޔ0,S���󧇳Ϟ�ᒨ�-��}�!6��Jyv�醊�^_�(�H�(y^����o#����X��3-�k\8�M�T�"`R�DF6ȕ� �,5�;Ҭ C�k���1\������k�t־9�}���� ���QHF��"��t�9 ?��{E_�7��!����]k�j*�Q��~�=�0z����o<���_TC?�];iW��M�cRii��6�t�O9_�v�(����ɲ�Y��\��i�,�i�W����7ۅ�2@�xd��,�)�O��
m�Rf�_0���6UT������1����L!��Vr-3PG���S��B�K_~jC�����ԫc����	ѩ{��X	v�r�9p��R1>1Ũ�SN�o�.��Vϳ��h#���`���Œ$��Agq�e.�K:����.���i޸�ѓ�߻�^�H��J<{��z@�8���`ԍ���fS�b-c��)�`l6M��5)�I�nuHJs)���N��ˆ�$�:�'Ǆ�>T�V�&͊e����D�.5@�'ɀ�[���2�) �d��@�ClѶ�PzEX�MX��!��.��E7�@<��$Ό�GAѧ�O�D����jm__Ů�Z�s88`�s��qgF���MT�E��B?��b�)�2�Ca�bM�W_���o���"���Y��
7�Ma��R��'w�(�"�@�/�|ؒr��C�w\%/��|7�U�J_�5�d �/�����/������C�!)��+�5U&�ĵ
/ �ƒ��EJ�V6zA���h��~6g�*��U���l�0U4Ep v!՚�K�F��H�VQ}�Mm�5d�3a`��J���'�4S�c���M��o���w;YF�����г�&Z��;I�T�|���Z�`9��v����f٤�
I�5�������6�y�,f߰H��������J�&�Ga��س��w�s��ɳ+���~���G&w�(�I���]�i���2��r����t�O���$V�N��.�q�hٚ3�!jc������I�#*�n�Puѽ�)�1����o��%ī6w����tvF�J� ������SYT� ̮X9'�䵡�P�0:�6�|*�}F�F�7P�|��5DO81�Ӈ�O����K���	���y�L䑔����5^C\u����V��v)v�,M˔��u��a8/�~�a�>�~c�fy����n5"��ddp�HV��ʳ�O��ؕ ar (�|�������}"~{��\��y���"��v�;4�g�l/������]#�ǥy���vP��G��������g�)���{���(�̧���g`R��,�uw(;Eޤ��S9�=�[p��畃����\��⟍�Qa�� �Ŀ%JQԤ������+��_#t���z,{�=�}�6!��j��`��5fg����������c2��`F.�v�4p�E��9��[;�A`��9s_L���#�'|�M9K��ϕ(�RKH|#+H�N�BdD�O�qO���H��gZb	DZ����*� ��D�X���ho���2���_��c y����\)ĕ.�`�o�U]�$��E�B�锋m ��=�i�sue�Es�ٲ���&I^L�a�q78YM�f�;U�NDn2#����jhݒ�i�_�w��O�t+)�N<Qc�\<Vu���*`!%���H"? ���̵���'�1�0YYu��Cқ�p��*�-����8V�!|f�x������f���`P�_6��J�ᕪ��U̜\��x��/���40Qe����n��bg�}��liɜ��ck��<X�<�MɧЋ/V������7�;A�=f��sFN�Eݘ�Ne�3��}�Ϛ�*'T.н��~���_�kq,5����83i�r�[!,�5�V�U