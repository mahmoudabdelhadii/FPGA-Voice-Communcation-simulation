��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��,�y�}�ǰ�=4d�H���`I"��W�`r���T:tB�T4D�m�)�	1��I�t��
��8(�8t>s)ו�."[�漆���]�~�]��;�O(1#5���D���d3�q	��9/�I�w`W?ދ�S"K7��5�,l��C���
@E=D��!
����荾Z�V�h��c,Dt��&�����]4w9K_9O�=l�uE�w����[R�\�zÚ�-J�$����åCj�[�
����T=���K���h�����,������#�z~��?�G���B�~֨1)��k��yq�$/ju�YA9��SX�{@��mWt������w�F��r���������O)�mC�&�����$��^_��|�����=������A���_"�s���50��-�ݡ��kVE~�cu��'Ah%�����v2ݲK:|�g���7/��=Q�u�~��qC���
qSa�a�n�m(�]�h-�FK�]�Z<��K�b�s��'�����C$Yכֿ��h|�[@lXJ�*Qm?�аR��(�v�vlr�j)ڦ��0p�s�bv��jy�-����(��N�vהS��Y�n)!��\|9��;#�o:�#��9|TWL��L2=�'���$ƫ���19�?�:H�A���T秧���,rJ$�p}�a�ڡ�rn#9���~�1e�[e���!������{�T�7���O�z�������쉎�<o�j��D�7��lS�ƃ���F�V�:¦?�,�:4I~P�o6����2
�ԫ�#��G롔�qH���'> x������>I�nN1.�yφ�V�ǹW�)��	�3���k��c�Rw�buRA�8����\��L+p�����U�|4�}��3w���n��B�2�Y��Bر�An;|ܿM�MT�[�=��Kv^��L�`.���kS� z@���Y�'j����@ڑ�Z��1\֜;���z{�ړO_�C��m��UW�˯�1\���-�P�DE��`���_Z��6��c���꺣���ĩ��6(�Rϖ���~]��\Yx��8u1�̪5�~߆!�g�T��nໍ!%���!͋��A�ɏ�ɠ�!��!�6�Kh�	p۝���wچУ@�,�Y^/%"f��ݠ "����i�����V��i�s�E- e#�nv�vB� �	�8/F���m�Q�ʣc����d�j���:D�&���7��oB�DTMi�@l>!1���I�$�!�s����y@��0l���ԩӌ�[�{��V�cr�䶀�����x�3��	9�f�����hpL���Y�Q�1GJ&�PH����8t��,��� OWW(�9@���YfC�i�9Q'�e�,���?=*!tQ�a���q+�+5�-8���K/ڢvŕ���|]DD�se�pB^V[���i��Ͳ����:k�"5�U!RCzWX`&0����~D�	�$?�V@���R0����װ��W�[��1���3kqZ0��>(fc[���iNbZ=q'{�q1$��_~ڐ�����9��֐�R'L�>���)�E��!�H9�P�W��h���r��ʙe� ��x���K���A��"
��������j`�%=މ$t�rm�DQ��dI��!�Pl�ި�����X���0E���̉�P����$�%�մ�*ާ�{�#�V����/߼�+ȥM��F�727D��|8�|���g�UJ��}�p]���G~�v����ol�� ��H:}�jpY{e+S�'� Y��j.C3U��(�|)��Jc�U�@`�[U���~gU��������-�1�1�,)#V0�sH	�9Y���e���"ө�EQ9N�h������SΪ�#C; �PY��(�7���8�O<7�Kiq�
t�g��E(��p'<qu�nI���1(�>���=�I��� @��{��*�AK_	rc%'8g1GƘ-��v�=�|\��a����*a�ۋ9�����8} �@qՈ��=[�0B������}f��o�(��PU�iT�4����z'+��Y������CD�ш�R�j��BF��w�����8�	ls(� ��sI|mC������w e���?yM�K�eڡ�1�L���\,����:ua�������R�����z�Nl-�1�mE�!_K�/��	ӂ�0�X���3�F�E���u2[�ɉ��(�s�X��7N�F��|�����{5��%\q��?�Ӄ=����f��À�T�O�/G@n��!��2���&��"<�J����2��Tϫ/PN�"�P2A�Ky�0���NOL���m���t���-ThJV!l¬V�R�j~:���Ҷ�!i�� p#H-ι~��M��GT��Ig��NI�qg��W���.���%�>M�y@���eL���j�э�^|A7��|�}�O�;��b�x�ʄ)��Y�H��
�di�hnp`��qsE_�PS����m��U���X���E5��)OF:PO5Ł�2�`��kv����A\~<6'?/;&)�������7�W
EO �4��qQ��G#0��KX��V��L��[����o���$s/?��#���GL��'F��f=���{���fB~�m���Q��!�T���Oh��z�|��
A>��k����� ��H/��L�ى�@�Sk�����00'�]�\k�+ll4�@-�3G���ў�/xz!�KǨ72��뜩�����bm�W�p��T�!�M�k��6�T�@��.��L1.�����)�^
����<I�%�8g�	���qW��P�|��A�>o ��L�L	��PQ��SKr?KT`
�� ���3Go�9J"��$�	�D��G��P<�]�FDZ��&�ʠ���+��� `��L��ǎ/h���{t4��I��4�V���ĸN
�����Yx��?`���-v6�'�Z�ϑ�:Ʀ�+�z��3��r�N)$x�ss{t����gM3�b�D���g�{f��d�'m��R?��?h��#*��-%��Tj&��lߤ����υ����o�}����n�9�o���8o-�6�Ve�%��5�RK�S=x�aGT�z��
P��&��T�L�L�P�/о�bs2�)a:��s� �w]�����7��3����N���p���g<ɋr��B�9	9�� �%�PW�v�{��D��,�s�T��z�������cL����K{�+�ŕש&����	��"T*��	��N*e��'�x�	%��63�׏?��G[y�V�>�]b��u���E�����
0|�%����w�c�ʭ�����t(��;��Y�"[��+���?����0=��sзI��腰��9T�6�u_x�^'��
����9��w��^�J��\��wIF0��\V�J����ѴҊg��O�(;���#���2��E��b���0��8wӓ�F��6O�:x��`N:/�v	K�Vܠܾ�+,SA�Zy#0��'��9�3�w뀝E���E�_���"Nd\k���7�@�����N��fռX����N��-��w*gb�(�ͩM]��C��[���ۛ��/�~��$y��~i��}=��<�k��g��Q�\�p6k���p�<mW�('SV�{@�3\���vMbK.]8nF�bDWx��1����
�SMX`Q���)�a,eA[�Ix��T~����������ϥ�EU�<������y �F�%��{a�UƟ"uH۠�!Gxf�B�@.��CXeO���aM����a$���]G�T�f���V8��+���F}@��\�'{�Q�l�� �1cU��fY.Y�p��!�q���<�͇(a��h{@����P�c����7��Uk�
�*����dH�<^IR�}�*�� ��6��Kë��,����G�����+"���ְ�胥�ތ�T�>K+ c���x�m/��	�&V�����X}]����/�z��?�p����I���E��
�H�-��nA��b�yE�8RU�|N�}��+V��?��-�C�������ș=�^g�Ҩ�Y�&�q$O���VN��3Ǣ���9O��t#-g���*^,��^o�3�'�,D�$N�B��y������F������jS,�;�����U�䍸s؏U{�ңQ3f��-X{�
��Dܱ!0��3O�bWe�3^�.�q����!s�`�X���tW�6A���kg/��o`��`<�~�\����I�@��"gnw�w����91ns҂�~y��b�/��l���m�� �9⁠RU��v�Uޑ�om��b��^�!|� ��ճ|��0��g� z<��ʎn�k&�)�h��L�a-���a���!�wW���l i�R��.г N��>�d�{��CD&	__02�!^���!B����Ҁ2ճ'�%�B�Ӕ!;M�k>��y��O��,��}�y�>�p�;�YVⲄ6*�.�BN�*�����G]�3|=�9��p��jH�/˴���x�y�-A�IbnI�X�{SX�j���U����z)�ydpXA�P���,��B��6���RN����w^ԫ��C͎4�R�VZ'���z�5q�:R9���1���[��w�)��`MZ0�q���d�7#QV�އ�܃e��,U�*l�d��FChD���ϣ�#/�E��z�#3�A���Z|��֠��VM�3�d��O�NLA��v��':���x�b��6���+7�"���B�����S�ƏZ����۩�V�J@���K�G�������8L�k�UOzu������u_����7 ]Eo�1�XU�	��oܠP�N���-��9̺��½�f�S���s	��0ܸt�z"^eu�F�� ��p��J����8m-گΣ]���%������*3��l�~O�f���e���#i_ Q�ONc^��Er�c����[�'YS�#h�LIl�ȯ�K|HL��U�ڲV��_I��JV���Z塦Bl7}�G�{(O��L�/�Ϫ����6�dV�}����N�ƍ%y���X��Ty8%�~Lm��wJy��� �$!,�(<@��/A1��0�BcY0�[�"�5���FU�XƔ �����:� �=� MZ��X��1�9���@���ی8o4#��SaϜyx�7T�1�P1h��h�p������͆������Si�){����%e���ɽq��ƹ&�{�a��������M�|���|* ���xX`����j&�IB�i`���� ���t�zר�U�4=_L	.f�x��p9ek���^:<���AJ���
���զ6�K�%S���s��e ��-Y���7�Yi��;hut�ܬj��e��:�Pa�/b5��DB9����rfp���Zõ��Q�Uk������H)��޲QO��[*?����A�R8$�a��;���d�8���{�&�h�hv��̼u�Zӷ��,E�_�a�tlSh��?����&O�$������`��=���{��¦%�@�됭�cY��5a��{I6��SS��"�BW�8s@nv�����<b�R^m�z��"/nK�s7;�B��K��	�U�|�� ��v��q^��2b����u	� ےAh�_��{�nb*_j�x���sZ�X�LS��Z����7q�l^���Ҩ��~���	J�[�Q�)>�{�-�F �1F�١ghJd@��׬�ڽK��3�+�lK�X6��:��f�6�������#&����ӝjO%��X�K��m����j�E��ӄJ`C����S��*�Qn��ЎZ8l �ԧ޺�<h�\.&O,���+�Q�YC"^g3�C�>�E���9�7�i\i3����,>�(����8=@
	K�!� +����N̾_�3��q��_`���X,mo,c���|���{.�k��@2�z7�,BG��_�L��984TK?��Cd�A��֢�r�`���'�������/Ջ�r%c�$��e�������%��SD�X�ܿ J��u�	�Bi��:�$�0ںनco/���ۈ��׃��,T�)�=�Kܲz�+=�.a|�L��fڂ�
��ԋO�۽����2��k��'o?��"(�μ*�uwn�z��)�L�`�gO�&����X�~��7	����;T��R�¡K0���>���t����C;��`:У�e�z��NV�p^��rD�<�X��P�#��,ߣM k]w�ݳs����ɑ����2
��9*�F���\
q�ƭ6M��ͺ�C���|�;��Pu���f\��9�p+��.Q����|
W��f0��g��<[�g�쎋���y�=��ǋKޝ�	'y$�v��4]]�)�CԮ�U�����@\��!�X�%��UX$�d�[�r�^U*D�>��%��3��3�zX"c�5\	�^C�����26�	��h����(էQ �!|��͹uLr�Y0{g ��ח�Q�������A��vm�c��H~��8IXXU��8���(�peL�1݈|�c�zx��S�Z���t��{oߔBk��e�_�L�V�I��":v�e=�#���M~)6�E���o"=A�S0#��g�`����ȱ�i�����*GE��K���E��[���=L	�F{#����7*�Χ�Q�]���E��k��k}Y�N�D�D�{�ӊ���`�`N����>(�}�{�������b�L�<a�Fv�f,�!��^Mq��Q��(��j�O��-J��-����Y�%&�2���g/7nC'��u�hƳ�����u��%�����Ք�Kx��H�{`Y�;(>�_)��7_-��`2���C�����qe;�/[[' �]�/� K[&������&�)�>��jHM���5@ع�>�_0B�%��dV}p�3G�N�+כ���N�ȉN���&�){	�6�C �r�P�ژ
���T٢������F���L�Ģ�p����i�v��b�]��4F�\�:z6Z�!��Z�g�{R��r���/a728����r@BOK�jB=�C��| ~G2��7��5����8<�6~���T�B��?_2e���d���FA�)F���=	͉ڶ���F�R2��T��>ݣ�ϻ5mY~ �챰�l� �@d���&���Ga-��<�e��~�����(-|��ˤ�;�L������2^���͗���d�Y(mך��!��T0�wqx�����ح�3Ų�KC/�!��w� pƷލMZo�!.�(XkҨ������A@�oZ�o#�2y}�BbC��eo!����U�}�>�����S3E��QڝD�u%	��ˈy}(6�������,L�Mg��N$���&�`&�
iv�*bNϞ`��7>2�3H��J4#@>Y^���u�|7E6�+o(4U{Cɛ��bjȇ��J2�Cb��,�1Z���; ��`I�ĘqI`���5^ia7�3��2Bx��0�,N�(F�VIΥ��d��4����̅��k_�t!m`@`�)f	B��nHD!]l���dX�QMh~�'7��w-�pPZk�& �i�eٵz�]���T����4ڊv�e�߻+�T�AL
N�/&⪠�;�p�� (xɮ��pY�D��e�b#M!�S�OYU�P�ˢ��9���41�&�%	N9��s�7���S~�]��6XU&�ʠ����;��qC]p/�_�L�t-� �¹S^Z(bt�뿨 �7::�-D+l�̂Y�l�C�����K$D�~�w�\����)�<���P &+B$	���L0h*\(xVhzE ����/c�<Sv3�MstAo��ͯ�y~A����7�@,*>iG삜2��CD��ĉܕo��X0�JHT�_����Hӷ0YK�]�Ե��@E/�h)����*�uLm��(��%�T�8C-o.�6`���]Q'2"�lI��5 ҆�Q�{��<5V .�Qإ-� ����⡅8j
�8�E9#+�Ԯ�89�9+���(b��BL�.A@���XU�����ݿ����`���b�lAx�U�t����;�E�g���-d�v���N���w�4�F�v,#ɳȮ�+�P܍�I΂��w&���{�����B�"VH�/��{��H4B���n�pc�ۯ�R3p�>�Î�+#6kA����ƅ�y��`a2mY�mh�n# 8�q��Po�\�e./Ay���B��w*�
2["��d�}d���!w���w��v�I�G��CѾ�|2��"�N�HH�����9oD�F�W�z����=-����b?#�巔r� #����!���г<�3�۾i�k�-6��+JI�f)&�J球'�Y��w���3�3�@�-y��!`OQ3I�^��ZV�?_�Ź�#�q��l��W����T���)�<%�<�9��Y�l"�[��&Yi�aG�/��@O��h��`@o3�x���t�|1�����u}�@�0����3�����E���W^i��zja�@�iR��-����#1�ѥj5�>4�e��]��j��#v�Sb�α�2�j�^�����$�F���<�HM<֣KG��n~��TZlH��0N��Ax�l�б�T2��1a����;���lPL����Y�Z�L�(7X��ަ�yc�2e���xq/��vK��B������q��>S��� ��+c�`e�+���T��� ��'Vh�H)��+e�H�8���C�KY���54W�r��(CJ%�9��oG�N$�S�\Y��
��
�-�:jG�V�5������}���b�t�zyD��VV��'ڄ�Ğ}���Tx�����i�s�� �;s�E��
�T�`�U.P���!��ĸ���
�B�8��q��)��;(1_Ν��EJO���G�៯��`�}Ua�Im���>�V�t��U�q.�uܡ��Yڥ�.�����I�� ��WBٰ6-����b�YA|�[�[���z�y CytC/��0>�\p�i�.g����7i��{'��[̿��UG�DGY��w<�)�ǒi�@,�E�? >A��;%7��Y����k�_��V6�F$ë��.h��%9��w��3>^���A�ʼ��z��ia�ER��"��5�jӘ�/L��=	-t��6��.4��Ѡ�$�\�1��N�ɼ�u��2����Q�ٴ�����
F<ax�x.�_���&��Z;ft遻_I�@'�fRu�ܜq3<���f�I�{]������<h���B)�CJ9���Pdh�q���K�G04�Ԟ�����q������dLd%X�yP/�.J�\qj{]�2��=�v+���v(l2#�}X���t����z�[�7q�_.��c�M���q�y 4�]lg�Z��rs��|�֩%Xw�Ћr��V��oq.j�ɍ�0��n��ES�ծ~F�xD�^��cZ�r���"��ת�Ze'q��J�V}O \zF���͈���_pJf�C���9����� P��{�0�/Jg����% jU�lL:�\�|���*�6�2���*�g���|�OQ�!jYt�B9��h�I�B�n��v�pG-՚xK��U�+H�yU ��z��
R(h���Dȋ�~GJ�S��i.*��ArOF���t"{Q�S�eMђ����IUe�wKC�BmE���>���^s�o�[\��,��j�BD��8o�K��Y�+��+w^RU{�wD����7ұsp/������n�	��xe?7�q�{����>��2�"g���8 Z�����y80��h�j�#���B�e�v����~�7;�Yu�˧�7(Ī�g��E�% ��4��gO���#��l�>i`T)|���2�[S{(>�e�u��$����u�QY��4��v`>�8����4��.W�2�S=r��}�]ڨ����%h,�
S����xk���Z���>�rF%�yJ�M�2y��T7�Y#5#� �yL��T��sʤ���K��(ҥ�DU��]P�-�P2�a?.�L�|H�7,k��+�40P�B1��Y��hK�ڠ���4!��A�`���nw�׀��Y9F�ŧ�h�*��(�}��G\��gj^�O��7��4�t��͸�p?���z�W�r���dU�(�W���\23al�9E-�e ��T�2���w��>JLD�=pid�6V}a��d����%��x�:��3��Wh����o`ayŭϹ����%�'�J �V?�ѷ���r�]��+�;�[;s���S��V^a��G�� 
��ys1��	���խH;���p֦�|jJ�����Q�<cgH� �s
o��V�|�{©-�C���a^A���s���v��~�^����A��S����	+Us���q�i��uǴ���>�g��a3��"s�2�!��z�UZ�a��L ��+����cdm|qăo�66b� �:��ʬ`"�i�:�i%*j^���F��W�JO�S��	ܖMȡ��'��[B;�>!������ N�(��~1�����ƕr��|�ӵ#v��.���e�A�aڵ�����������2G�������'����_�!�jr@�q�����x�R+ol�����9_�ܝi�Yu�1�_��U/8�I��N�pC�ec��\�O��ƣ/�/����ko��_��%�x�.X�Q}L�s��`��x$�b��ii�سUt��7HrXm��D{b�Lh�P�	,���������qd�E��m�V���h�Xb�F�qR.�s� LW�!v��W�}XT��g��H�-z����a.���������q�n܍~J�j(����4��~g�t<�-�b�W��uRՃ5`�z�kQM�Z���u!�-��xhH�Y��Y)����O[�Ԏ�f?pYA<��ͼU��Y�Ě�T��]��p/Fg�/���I����	Y�aEi��ӎ�|��*ڄ"f]О)fR��,$��[y0DOT��)���R��������;e���fm��6%=��S�oi)ށ��(j�5��`��r��)�p⋠�P�Wz[k�q[��y��b�鷺�1֜�v/�%R��{���ɔ��x%i������
��'�5?��.}���_^�?��l	�R�C)d���Jc�����z�]��e�;pƬ7%Mo2�#j5�R�apt�HL!K��Ve/j����
WL�0]�� K�׼�m�Mw�ʣ?��8��Gim�n53�2�q;5��z��`���=H ��V�)�1��U��)�p����d�Y�;���euk�}�jW�ߓn�E)�\���<���QFI'�tK��ţ���;>'|({��"����m��|��
�����G���o��� �0%�g����%Y/Z���8]�E�4q_� !��{(��k$4����[A���m]e��,��"��=�qM���2T�}L~Ttz�g�<�@P�?{���l�/N0�Hr_w4D�cV��D�M��Hʃ�d��e$򇵛<�}
h�ԷCo8��;q��PS�����x���<V��<d�I��ǖ/��:B4՝ߓ-� �|l��s� zU>@1�q�gԣ�<y���1o|]rຢ�!��,��_,���X�Z;V�9�!�hU�n��<��0��45�'l���&�����9}��*^9OyK3����ER�W�OR#���ͭ�+��2��6�dv�ziUe�Ԓv|XW5���9�sWjN�r �z�!�F��pȘ�yZ���Q1�v�dt�١�W�ZL���ǾTPY�	��B��'�$��s�C�jnJa��z��6�	�m��25KB|���0ҋ�R�K�ׯ����������.�������yc�l�i�""`��GCs3�eػ�ԯ��lp��}�1��.ˍH�E7�h��O�ʕQ
��(8E@�'��:-�	��v�~X�"K۪����C<	#���©�.y�t*!1���yHKj0d�ߔ����"86i�a�<&�����c�Z��	��9��2�W{���,�A�O�l^V�ӷ�"�0/�	�h<�D�,;}��E�m]M"4ѦT�L�{d�."0�F�9r�\,�[:
^|��	�5+�,�!����Õ~gk�VglT���v�D8N��);W[e/�Y�5��`_^��=��&bS���f��G�wS��WD�prDGwQ�+��"�5BX�k���^�'�<�����M�*�������w�2�)���Ar�����4�hp0�v�V��C�q7�v��R�f��V؆�7�R�"7.�w_�a�zL��JZ�0x�2�S�oX��C��9��(��<D*���8�Le�:&�?�h#�t2�(���",<�uϟ5�l�T~f˗�{���E־,!���n.���_'/\TVx$X3�&a=�n����M\哯�ɢD[�lf�������P�:z�is�ʠL>m��w�YB���l��0$�+VlחE���Ĥ�~��g#�B眴Q�L.$Q��B���X�vk���d�WL^6ʄR/����W�E�pm�edL�`Fx��i��Kk`�{����n���������E�n6�$�Y��5xu�����NTϫ7�s��6J�*�آ�*1��F�W+oY&�%��ʀ�ͥ��!�����3�8���F'B)�N��5�Z��s{@)k�I`6�uci�c�� �ZO�o����q��ͱ�u��:ue�X��)��7C�m(l�?� �\�yB���.���5��Xǻ��;^T���ȼ⛲Bm���q|M�N�Me�K%�[X�x� �hi=�����7}dtkc��o���A�o����t���wp�%MoV�υS����.c����"U���.�!�1&\q�xVG�c����
����IO��/a�c�''��m,�r"��F����;zூ��}����;�P9�G梕%u�٦������jI7IQ���X�BYF}�1�G� �(���4�1��(�EG�q�yILĆO�ƽ�T0�/!�{�h�T��.r�0����u��W�מ��W���r.�I�̑�:.�]=�����Z:S�׵���.��7>�"�&!���U���βM	��Q�&�XV\dsЦ��F4-v�t���-.14��Eڨ�,��Y��N�"��*k�8+��]����.�o�(Z=�/V�w�L�\i�/~����y �e�bgmrl�����w�}rZ��X�g0����E<��0���҃c�,�̫m�XYտ�J�Pt`��C0��Y�����g���۫���Z�
�2�l��F�}QTI9�Q1�
ue1��b~����~�p	�q��!�ٕ�`���G3�h�S�%�d�va�.A}��w�.��褢�W�;������������؅s%���͹�+��m�%�+�bGA�0�@t��h�";�}��1H��l^���1�7����+Ǩ�P�޺��鮜�r�D�1�^�"���躾@��4?A&�*bR�{,� �{LH���;����$�(�3������w�Na��Hp�^����{��7h�gQE'f�����2)h��D(�������cyc8<@�d��cq1�݋�!��@h�C3}P�(�QT��743�-�@!@+|��D~�rjܱ�96��BF�h�۝�����N���2�p�,\,z��C���p{do2����,����3)btge��pď��U�W�I���Q]N��EV	�/�k��ɤ���?��l$�%e��#k�b���Q���0K�U�׸��D�É�|�n��	�9a�k���c$K��W�}ҷ�����֫����z�I1�]	[�^U���i.��7\��,i ]�Lcx��+w�5���=�^H�sz+��;)�x�0�y�>�����n�!�z)
�mw���M��B�U�PO���a���jw�#�^�b�Vђ��?��߫��`���r�H&�~^�Asr�/1��l�6wt#��n׮@�(ާ��~���
��5p��;�eB�-�_�2���h0օ��6H�:��q��|g�����C�C������9
t7J��ݖ��v$��X�=����]]++�����%��l�C� �ܪ��w����&?�����{ҙ�s�o�����[5:g�ܕE���'�TD�c7�f��d4��7�4�Rj��t&3�~�p�i"��r=�r�<ՕU+ۿ�?L����j�gsg씆��v��$�!֎�#�P6���E�[pT}mn��c���y>��A*�
�Ƕ���Qҿ��2���P��6:r�:��e����"�U�ߙ�f�,��f5����mJ�Y���I�U0<I��@&ݥ)|�e��8-������T�8h%��$9�4�Z��6ڰ$�+��*�6�.!.�)�h
ʭ��
��u�`Yh I)ף�ث��Z��k [�+j��#�)*��/���D��7�o�*Ɠ��V�'��p�����2۰W�R�&^����� 7��ƃM�,<Ӟ��*;���� ���؝���qAo�(C[��պ�X�<U�դk�D�
����pJ�+�Z��j��<�Yk�L�f�~���ַJMQ��p�B�