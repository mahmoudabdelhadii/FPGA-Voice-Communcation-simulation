-- (C) 2001-2016 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
KgReIeriBJW9JzZ6c0Sj5F6i0p2zH7Il0orVlhLVI9cVkafe/1m1BjwdBCp+mIQUmVoVAi/Y5rnh
R+/peeVUxHjZeQi0CO+1jtvKMCFcCpO1bmQmv3yLPQuMzjTqFnD0kbVGu1dCNiJvItQsWLLhA3JX
XJ4PSe9QGhr97uPtUwLBC/FXJG4H1PjF0hMwZSaEhNRETQ0UanYhCbZO4jVBlvnf8Y4xwfJpzQk3
HQsth+3DJngd6AKHsoph7P0Uj2JxW30pT+cInsFOh0Hsg4HDoz8rqgnb9/d6ehLX9fxGrpYQEVcP
W0Fb3WEjHh0zrkfLLsicm0hX63KUqzPUIq44Sg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 3840)
`protect data_block
pyg2UZSvlChfsS5741nz0aO3z9+gn7+kS+X9o7DgX9QbNlog22Ak3ViSFhXH7I0pflC8NRnJ/OqA
WRjj/krsunjPIPy2fzTUxxpBK9Os6vWa1vjaWLntFnVh5bIrUwvXRxdjxvUDZvbHJasfmnwpuTm+
WvGoLknWCi0WG+hrNbpkxOucfGsIsYAdvDXAqIsG6BElexag/UeAOtOWmR/QbDZmpRdsC0Y9vQTk
ypbXHWdVBPd8EkBAB+WeMiAHTZUyy69l4CGiyVm2CXPyZYQlo71BEX6TOMTLZYuY+kQhRwhwlha6
WnY5nlJGbRxgnrp8/y4oe/vxLz8thJ9VI1UyGZgJElyCxgTeahXrj8H6ZzCK4H4JH6yvDUFV+ML3
UohDLm2UBaJfICAWoPRkIBXcPZ2ucA8xo+Q3HwFRxUXXSDnRBBzn5DchyFWT2965mPbMPCoPAsU8
vKS5IeCxEVW2C3lIJJlFX1nlw1M476riaMIE6af/fSgPhKWYxMyWYJJ/vJLE2RxvDu3D9L+YcwhN
AK1jn7VXn+veF01TOiM6b9XP2ww+uMzXS3G+SsViGpNLTGyigS3jIw3NqowP+WMXpo5in5+z8ROR
IrERf6Me8CKUh78eZG3HEMFy2iBSOY84v5Qv4IGbb/F/xTWDCBRvW96yJQgYH5rG7uGEQ0zzaUX+
ymlNwWgD6dW3r7yuDmSIbj8LL9tEVzMWp4TjlaEE9nULr6EkK7lJdprF9+W4Q7ftAUfqGo21cVpO
M++EPtBtcEum+VRyWXQDH+PFB7+H/kSfS5B3IAucE0XHRMTeb4Q8yGjZkbGp6w6kI5pR4MOUxduT
SiPslP5sUI2yL4qFfjw2OAdnhGrTTZ4z5HK7lpCcHUdQvWwL60NbRARKaQHrJ64GPmAXhIjFWp4C
wAM2y0qR307chhlXk66/x5pbrwxf6VzEKgJ2TyDdzSeZwL3Sww3XtIY7ocVtZ4TkNhWRD7LPwH/v
nOzQmKgAl7o+KCT6Taioc/PgVxcASbCPXRCwYncUl74pr8dycgjPssBlx/gMFee5gQ3vMlc5iu14
0O4nZd6aFHMjUCUi4/5pV0ig3BSqvHd3r9VNHWthIFNjUSIXmVynEVMf8lxqkDqJjoCRZLFDZKOq
ncTdpRnhoXhqG63CFOsIxk9cjxEJ7vCeMcRL1fAofId7+WXU8CHCOkWXTQzOr0KzGUfD1JOf1e4k
/62psJlA6D5bgJQY6ll8a033jCtfQmXe3SbPUQklSrBAxryXYoXN89z/LnFiAUzYrjliEvwpC316
1rXEnyusck8R/kF+M43mNBWTZ+TEqD6ouI75ygvnGbKT0YJMXEcrqK5n18Ec6icYU5gFcirJZurm
5yoYhOQlWxk7AlXgWCHRvVR9QAfyLl1W43NQhfdZXZS56KniN3AhpnKju/O8PpqxCaE2ixHsCA6j
AJoOZR1KtnzPRxO+3Pd2WsvqLd2mXUYnj377erXYKQSZO5ybU4pVp51kjNWQpkpFH5f0KMQ//IGo
W5KFzPvlSRK0Td/3BV4g3JNQpILl51lGs7acfOObMNjd/YJodpijghX+L9sQU7PwWu6k2umF82zV
1ygO1MYtxiwjd4WSm6EmJtfDiMJXzuUlEgsL2oYOpgrnAWPEZETv4lEIRsoVx92A/Buc0SnLNbVb
8ZQYdlffnIf6ubjiE31KqvSaA+A86zu8SBdu9YdB9z74PWmuW07M8aruQvcYveNabsZF/osGGUt4
imOjbuLib6nELpooQ4cgTSkq9NDC+BT8EWkMEJ9QX+oa8VWIw7NCfGmTNbFmg0liMAta7tZep4sH
dukBAJ9vqTubbsoS+1Ajynm47ZRCIYp4b5uZmlH220+ae7eXurKh7AUbbQZdE9m8/7GVgbRkYvoD
mP3I4z2UN/RuZi1/nHHE6WeTZLnDR14Wm8+8TbCJ/r+UU9welAEvRS+UF0p9t4puXAVFS3tSb9vv
xp0tugvXrR+5t4+3ahM/lvjFtR//7nxS79CRvDeifDJyRCi1ramcvQybgW1V43MeWRQI19EIz5rs
F47tj1PRMLrVOO+w2YHALaPMYP6WzOShOh5IvL7NDHkA0BVKX9UQ+e21tgiIXh5ZgOfLqVjKVet2
gNOyXBrXJSSrWNVJbp8OrpB5yqdzXBtxtEYAbbzGe/+VCZEVO1GzHVHPkrmkmjl3VjHJhHeNxG9m
Anf3ZBCcnK0NfEk285NzwpHS76ZFza9t/YPnVS3/sWuUgKv6ZnwmJL0U1jT4Bir+hlkAnYV4V5Cy
DUUBazkfLHh7V4FwxkqFge18a0W0YKd9BMNRsqG2zUFVbpyCD074tS+WZ/ViMkm2QLzaMMnynZM3
Y4aCVUsck0ch5dlmAtfG72yzeAwUEL0cSbNgDgU8RvwZytJ0Kaw0EFGLDrNYsmyiVcf19Jq58D14
FRVPf5kI8Lrsiu5jy8SEHcTtozue2ZHU/ktbbd8tCH/RXG9kl6QBNNUta9WCmmUOclMzAAk/Zn3m
s2j2ISUbsbrgy/8yvDBCJz8aHqLXZt8SatWKmYzizRBJQchHzf89ED+a1oHh7JxL+Zk78i92FVJu
cSmbnxPHRfdnMkc0NauYQ7dLFZR++4MuEDgho8+j1zdnwcIWo5Bwpqs9S82tZk5o612p5GAIbC9U
taz5zeMEMOGmVc4RUO4Zy7NPA2pbyOkvnFjPC7AXhRV93pQnq4dWpQ7vxlA2MyVMtj8RkHNr0+LB
OoIGnVCbB+hj0SbcuChNOh+i1gYUxYiYDNMwoF2TJRIBcUURsHe5XbZvrXoC8x7uhEuf5oNgDc63
HojQvWDsizLi8aHHPYLjUwqkWdSebmQKWcVG1tMdUgH0i7Wz9tyC7LBIjBGhVeyUmqu5hjsRDYaB
9KhBmYC/5XEa/dy47Lg3X/jT818RZESrfSY9wEgUi7DQvm1upbr8gIty7zv0SBP6OiXyK26m0AxM
cVFvQuh4HKTcrRp0EHuvEK8UX06ppqIVh/pA0X+4DOy3MQ37MSCtOAQkwjYSQ4B/0MpR9wJ9fSqx
YBq/lo7pRJj74cPFU08xfkHOAiHkbEC7426WJZ64+oNvhtlZXCrhz/0JxQA2LeDAjPjUYGUOnhCG
8GyEaBQNrt6da7VpNYKAj/heIHFs+wnv5y3bDk9oYyE2OQaATAG9xR3MIRCoDS1Sr5qfSRj4s6mr
7eZxkZZq7f0Ph8a0GDVO4sPfBdTg6RB6UkZA92EyI29E2FOxGa3MiA0bC2NfPa3cIvdtRdTXd0Qn
3MGsfInjKr/3KmU07ufPrMItjpxCab5h3xT3zqDayjx2kv8Ozqj7EYhlU4nxJOlrikOVLHQxzNc5
L4BQeVlF+e6l6d/UKQbcn0DXy5nnKxw5AgYBfw75p7EgtoaYwvpu2r1ZDyv8pjMteDWFMnphKDPt
q/kGzHIVj5fGCv0kpYBnmlQ1xwca4StMUibUZYQDfSncG0dZZeFnymtPyFp/II5HA8XhNMIe7NoL
Zp30wkO//v6n0Wvux1xdeOJ73/L8rkCN2v8SR6updg6BW7ia2hzkHtrCo5y+wYsK7DPSZSRFSaKW
ATWLosrFKSNLpZ6GHbh9g4KtIK/X8MZhI+vOQYTR+xbDhWiefShsIWfa6iaonVGa0RaQ3DGMofa4
LevBvsm09iFQ8LcMWKPt6N1deIwf/bR10GY+By73bWFwKFg4qO3dGykl5tpKWcT8mm6i3c2uQd6d
nHwdM3EpNOMii0A4xgODIuSWBp57n35SUt8ExYxArEh1lqP6ZEbi9CniNFipDf9HJW0jCP6e3oZe
76FW3skIxcJo+zqSEukWna/mjEp8Ymj8Cr1xq61g+61bKmY8U1aqXKug74IVfwVEBQ26NPnJTeA0
FMWB0jUlW9dczXizeV4IxB+PGwFV1XzdqQOtzm0G4T9Nks6EXuB3dWC9lDv12o80mIfn47gH0L5F
ZLse6lAKaSXb/z98SB9XsaEzYYjC2qIRKRyXRWvM821EbcyePAGSZiinNo/a2w84P9ygOQoWiifz
4u9TDkmvEkz4/Wkn2M0vcHQM800eHl/VJjSme2CQ/YuGM2qD/OtCZNlQpBVVD77yGonbbRyd8+Vh
B2HwML54S1OtymtYTqeup2TNeZgnIM1fy6HbaJWOCwLBAQquhIaYCM6cR9ZbNRV8lHWflrK1aH1r
tIRU+RKUV2PqHQHnSNWL3j6nR9spxJezBYrp5KGdjQJUZQzXhq/UsgaD8IkvUmL0RumG/O3/caEp
cYEbzSgO4SaZBQT5eMLO80BOQ081PBr9RJHVDTyvekzU5YxO35OLbo3R5qKPOyV1aIYSBTf66fre
snB1nXpZL3MqaKWczYivDF1xHV8VHMucVE3L/K5u7EcpqoZ7y6atHy2zyT9ocyc3fzJwKf1E5E0R
/C1v+m8L4losNtZn5Og0ggEuxqzClEgKGvj2L1YgFtktczpctosjgslBgyqZcd64rjCM7b8F68pb
3mZfK5N35aO0WPxU3w1C5ZD5xNMp1yfosm5sy3+I1GBVwumh71TQqAR8rV/uBGZIII6pNc9eK5Eh
gT4+aJQtamqeICZYdW/6SMTLOTaeZ/qk+ceMHMFo0rq+F+3skpLDR8efDJ9kWcsiAPLPfqkU0p5r
YRhntOctsUY41u66t6NOBi8KIHgA8zpFBqZqE+/XqlMX7uFVY2fhLaDhCfQxL4jViUp7WTf53M1T
ZIeqKf5WL3XVNvTqTRtbfSoCOj5E/mBp4aMyWVSZ1PaQXFnvkYqla7fHBB2Q/3MhRweK8RdsT1Y2
xBO7g1xlb/QREwp8MSHNUjRX+bx5V3SCdxfnjpqAjUhJzFkfCBjqgIn7PaHrWigwAcIvWFtQJ4IL
ji5oIQ/sAh/gCNcePf0faTHunBHFpeZJFoa09bJILdUXM5D9uGqgfqr4BmHvfUSa1hCJkHwW9iOG
7BBamcNEeVqhJN78pDqWEMClsOGS+W+sT1dEgEPY8b3a4rqgkRhuPTI22TPBbQGtXNWXjwPsCBN1
8ah3tKVxEEcp0C9e0NO6qQMte2+iQ8mSgPNbzohTomwoViNaU7ZSd+li8A1qQ7t5aAt+6NwMyNZQ
5OQY+GM3WAWSDZ9KrJ/ObcfGF7v9
`protect end_protected
