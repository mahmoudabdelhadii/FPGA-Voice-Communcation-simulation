-- (C) 2001-2016 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
Xi+IEpabdZLgB8Ct6x787M9kEMKfG7BCNbWyJk4qV2O3XWrXRdW88RYfAKbh2Yumvnmp6oZ7JZBd
hJEX1uU5VSFFRrmKRwP5sqUdxU1sk96Noe7TY6jlfYx4XiTVTvD0/ESQoJXvWiqLCbUX9sMq9iAO
X93fXQmTm5wfbTG4u/OiOjtDNq6870DuUQ6pWZWceNgCAw1FtNw5k4KpUMHXH1N7l/f/BM2sneDT
kn1E8qPRJL1+Pp6kF8shNVbUva4wziKFhSS78d+CjKxVWlYwgq2m2lwD5LQbmVHqqjbDPqgtE0ps
FMjmd7mzMXW08MzFVDnMXIlSiDS2cwbZ/kL+Eg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 5056)
`protect data_block
EUSMUFtpBjVdhJx74feaKQY32iZ++h4gJxOkMZgU7afUz54e1XaznK/mhwILMDwxEgK2VMqEn47I
P5ZM7WkGv6DfHBOyh5wiO8828IYw3Qrw2moRv1al9pU/0Cr4tNHfllzPOkooLgpCkr9iRYIRIOIG
xdIYpTvgY9U6/QgutZY7YmN/wr7kWj44QkEfrtt/UcTTL3JCdR2JAqjT1cwZgjawr/jcd3anrWig
pLUSrsU6SqUsxN43X8Kl67p0hNmIsoMh9xSiVIFVTEZzQNKSZm42YpfIeYjR5MGTIQaESwaAc/x5
SHPNNv4HRSpr2cTdlMbUDG02OPKgPn8nCDKooHnRHMGXaFlHRLdza4i9q4EFnUcb6gnmFfZO+tUm
QPrqQSFNUFhGPYNJpaS6HNABsx4Mlax873yu95vpHXrQvTJXtJ38UcHym5BdvOrf1JYXFfxJIdDM
/H3+77fZ3/NOQaROUHKuFEwkzNk5fIwrneMPzWopQ3ALG5OagD2TtTvV6G6v+QjDnKqA4De985Ws
gWnARLo1w+3b5HXwGiJE+Kjjrf6CRzN+3b3cjzpGG5nNRf47sM1Fg51+hg44x+2ZYUfM9eV3fKUY
VUoyArbZpTlLVKJFNjghE46kI1EWAUzrInxgH/nNPYaE5//Nxta48yi7tTDBGF0on9Rk3h/OH/9N
s3NmP7Mm3qXcLJE4XCYdk69dmwkbbPevoc5eI8FItVVz/YA4oPfJepv0IgTlOCufSDkyPteWueRX
DADcoLDNrIVCfg2dhuDm3yFRQE6ojzbJNlrULX8rliBI1n4e3ISmU31u20NTOcusEcXiMiB8sue6
UKi+urqHltQL8D9DKFyXbPtuQeVDYeFAYO0ExqznaqlJSmwgbLdDW0s63175AKb8pH07HZcW71nZ
VgXPPOSBPHq8l/M7U6WaMYt8EIBrukKFzNQYt/pqYqnPtTnFdO/UbutlxDGPuxfesZMT1oShSV7c
MjRe8oCH2jUpHKk5fZSTaVD24VjXZJpDxmprIOWY+slumhE9EWno+LDTzxiXNPFkQ6FOCZ6QwdRN
lCiSztqqGlzmrxdNh8jJi5UN0gj6c2CtlYBgxqEiSIFa+EkWzqCXe/+9fvDmckUEuwDcf0+V1LCU
dyHyKGvh2URSuIawgp8AL8V4jCTLGMItKFf2p0g8hhG3cEo4NTFfTrQUV+5vcOL8NiBECkjppn01
zjtpRoXy2bKCTrNq52oJDw1zscOhJq+JxJppD0La1JPVv2VLtij3G/bAZ8LZE4SeW/eIvMdTR1u7
gXF1gUf+8NqgAy3enpSuPpvc2Zys300gqsxIJaD563fhSfvo5/gGDN9KGZ4AghIsiDsZNhC3yi78
2+3QhhOgTmspavd6nF8VmQ08S0hNTSnPHHYAYeUXtAqwoZuBk52FYnrW/y5vk0ob63oCxQ7xm2AB
DLqkW7uJTSrE0rEmWOtVGy80TmU02zMbAc0ryu+w45TdzUfxNd+yBvSuuuKglTdabiQD7v7jmMv5
Qu4aenzXC1orTo+B5MfrUqS4sJyngf6FXLsw+w2aDU+w6ZDbJA3tmDcyJPVl34PQJsmICb+7EC+m
zoBGeIo1hyBNV4rtL+njQCLIwzqiXscaNytvBveQLG9rCEpCinr7v/pJvgWNs2owqIj4MCmnz9I4
H+t8avhR5gYxcRI+g9dqj947ye0my1Xc199fTF28Zy+b/KXHUaG+R6HPQn+5P1Zf/ZPery9KDlQs
O3XNerpG3ROQm/o6FH7JDujmKpEqYGK01kruNqr/kUVbQCb59OQ+ENIT8lsftUue43hT/p8xnsW9
xfUSV4YtiTxGUuKCP0njorJWBVXEE2RlSLZ7mHt61Ec0HZ4k6VogV6NebU8/cgu54Kh7nmt+nOKk
J1C+pJi9vNAbRH2l+sCkIRuzI7smvsEISEZBkjKcXgMDN4zN89sKqxNItjwsgZT+XnAn9u3UoMwN
vP+5cmpdJHN1l6EcQiNbeoLK+aG56JUf7JLgiIrlUPvspF7IwukobOfLwMr5lFFD7EZkpDW7dtSr
xWvXuTeRPI17NPMlBj6Y+2Uc40J+2c6evlKtxhe4CFNVLvKLNcxd+9NPHXM2qvNuGuS+z29MIYJh
+xkS7TXhYf3WR9pxlJCQhVG/FMFxqGOUAgwjLHh4ZYYLjYp2H1KEJxXo4bFETF8nR+4smRleOzxn
R3EbKL8/GHiFePct3KklgXgkU2gAot3E7NUugTWUZAk67HIs7BmulKJdgb6QDcpK0m7ANsktx+C6
MhpJDgd3PJJ6Ouaxplztr1WvXTuR14XXqj6hLmKhe2jyGPFMEC93xhXMwtq118QqxdIlE0RQUFR4
LDDMIo+GfkSybGgPxtqjnTBOxoRAMb3O/c4SnpDta+nkvjrnSjf7WpktW5n4IMau/6+Xp1JF3Jr8
6RrIJCnP9uPtOJasUURwlkvuMAe74eEfraEXNZqiIQQySFI5wDJJFimPtVyNYJiTi1ENHjEhj1TE
s0gHCsnV4rj9wa70LdUSvd95BuSEwaQ+TRa5FcJEzOiiVuQZRqfonx7fu6yYmApRCcszl9333zgB
MMhQFKjDyJA7noCBzc+AecowB+mCW7WddGUKEB2EpObK4Jj1fOd1cU3t2ZBn4GjYPna5SmiXIAex
PsxpaNocrUvd0s3tm+ETvLmy+GyEttStJzMk9VkHD40GFT6Q/sTMBlnXjG1PH0ojc/yw4onzavVY
R1q/5rtDuTzCIiW74sapZlCi+/iyt+1QQe9tOsy4ZOoPDcJGGNf+C3JCbEsCnnM7gkRFA8NPrnIE
d1EcF1jv7WmK3Kpu5h1eeyguN7alU7e160eKE4vPtTZVarQginQiCvtnx6wePsgqydDI1HIVRexG
azmJlIjBDRCUMlPm3CGtC1VBFC22NlGOKDgSrrYtcj9JHrHnMUEROvxI2Xjq3oJFbLvWbLHKsV+x
TL2XGuV6sZj6Hy2lHmL7Q7ezsHSYfvPPB9uQ0eSLVJ/RgfgzahhSGZBD6Z2ru+yRzy9e+R+dyLIw
UMHHGmtDGDioFqKt8ykD7UKXnIZLMxd2fxTTAXpOgTWglTnmfUUvjXxTlBJEW+d0yxg/LdRbwcsH
quvvqDpTB9++Hann0x2iXPTgmfhnDPqTlKt3XBkKjbDhxBsgTe1McOmiziCzmybdYHI6vYkj3VKb
1Z1up7bVdMmbcTb/6dRL8GNdOrPotqK1JUXJa3mJlUbenmxl9OM4rHdvh+qu534ml12NS5n8k2pX
LB8JVxrXuLDCHlFFyl++AkG1Hf4gSEQFHk9/tGVm+qcs5U5VQD843GbakDj1+rwn1XvRHXfrPaNy
ph9RjMCvZfPdIjVn4kvhJHbXRUkSpPglMBLxpZ6g9SlIiNCPob8iUP1n3Ur5WAnAuI2MA+wnYmcc
znhsbhvum3i9/kFrv106Lgz93SP7qWcBW2BruwU8+RTc+g6jAUpVJtbwMvV4s4iOumcpbEUxUCXj
B2JT39GfrRtV+hc705ShbCtKnXvP5dT6LPJ3Wv237ff7BKkcNjLHtAWrURWqKP/h3A98hV2UsWrw
r3vMAy9x2NL+HDmfxFBESN9y0tXmJpVCyOP9fnFP23s7/VuTrZ68egJ3K03ShXDhIlw/TXprtJhf
A3QybXQ5P+Fa5Tlpin2utRxkQ87QP6sXpMG2Qb7h7KgiUK8BhI5sZGWD16TJvoHD9xVw635nGMRU
xOqWRuwQk9CLkWDZXmPp31OyYZUhUVxjY2Ne8axm+ImoWHwkZCT16VINA1e33IU0OR6ZIjplkIbA
bHBll0pTWDSE86PQPg88D+nAeivTA/rgQnXzVdmTFLxggaFktZw8V10sZUParhxkY8/gW4axBckM
mLkGSjzQ/shTODaNU7cV0y3nWmJwxMZ07lwV5R/P3QbC7mRAH5HY/MNFXNvCZ46tDAla0k6vcOSh
XDFvLwlHWcZAPlb4LtPCEsrNyoH0H4nMEgb2rkSKnJZNLOJ3x2oowim12uO7063YTu+CT/6kt7HQ
N7VTl8Ds2S4Xm8U2HBmkO05ub+n32+u7E4RQe+tKC6jhYBfIcerREOoeuWQYh5G5KPNR2fiGtoDd
txrYNkyrVS/FUoyAu0oTDbN0xQPAyTdGqyaXCD/qakNnSjtVyLP6ltnF4HJxH/F5/7t2WTfK5BG7
W1fQsouBfHF2uWLLeWZpb7UhW1B8WnIeBk+CrbL5T8Y/hq51w/MuxFmSxEyesNmXll38yHuevQtx
Saq/H2ImSh1Eyn/re7Xg9Qzlq3nc2JaNQb98fK7GZ5o6fZ1VePyjoBb3fdXN3VbaYqj6nrigxLvo
bSTKkUYBnplcX1vScFLBQ8SQsciOQp3HYEdnQjnDjeduGaGdeMSjxqTn+hkzI4BEH6lj2rt8qWb1
v749mwEvqAB6baxhlzJ9qMCfwaN7Ldp3xVDxx9ZRCXmdJvpEvfpPJ4F0Vq+tz3DIpN2283QizQuY
kNCLN122QGq9tkc++BkJvuFEWhnpCq4DsuWis0ruecDg/w5I6F/NscyLc2EsvkF0N/SFAm/56s1R
L04w1NipKNHT1NJ54T6kyR4byC6nHJUzhPmRzzT3rsRx9S4wiSK028RYxrw6aDv5+SVYL6WPsoVz
PlOqveKyn0XQA/7qeR4LV4xRjTO4BJhiiNhSmZDE5GP0gyKKzVEWK6Yt59EK3q8stWseCbdQ3VCm
fiKqMFU9NqjYgs0dIsM8vg65+dTu1k2CfJjz+eRSpgpi/YPlmGFNg1/XZll/CcFGDzT7fNnFeqWA
wZ/oTxH5kqZV6/U+ApEfnyNnCLQVEGEaIII+KF4vfDYK1H45Nmcks5X2r3mH8me8u175sgd3gRYI
LOfD18s2i9xAJ+q7s21EWMJx5qtMwozBkD9U5JxivF3bQ00BxMHb02P+f1wXTTIgCM3CGOdA8UI4
GtvYybNqZFKlSZA8h4uPn0ZCTqXfo+Wm5GLeDuEKz7ttj1o8i0WvUxIuUwTpXAF9pOs+EyOkxtPA
aMlhKfXN2pl3j51bu4rsyPJHsy9swgbmJMfaKDZq+6oaqZ85lioXRfxcGc6J5qZGpH6ZJsh1QbXo
mmeifntX9uF9zszXyyVU+u8B6WbYqKa8L+s7+cDHIGZJQGyaISAfys4MtCQKvGtLow4Erf+dJ55A
pyyZ0kvQtZs33NiQuEJ5F7r8LsVZsj1liBzyPlXklXty1J3rIC507Mbkh1hEjuPTr3WYs5q1WDsS
s6jjICqi4LrnwSa4Mbgi9bDLplbYFslcu76Ouqfo17mlehBSkQ0SSDcMoEzcVUQdHP4DKO01B2eF
7lRynMlIx/aXl/dJ7toONFmOVluixaT665/5NSJzFkt72NDN7sDw499t1ffJNlv3yY+u+RhHTz4Q
NyfsdzIHRriBHXu4FQJeHWUqNOvUxemOl/CYfK+9e/s4o9O16dDeP1KMoj2NydC5swAcvQ6EsOOc
AVW6GvEpnE7OvdEqbS0Wae70MZM4gOyvW/QS0JZuv9eQJVGg59AjA5ZZAAJWQKJ5Foq2a8J8fwey
N+KAAvMhPoZyZ+Enyi4V1G5JwXREYNe6BGZ2qscZMd4eHNRWxJQZ6g0jRvr8t8LHuPi9laUuTp2s
mH27N7K8aPwZizwVlfa0ggY5k3tvm0zSFe+XwLrjSGF4bOF7+h7+ZraOIqrINDJ+MVFKyFrtRfjL
1csem0rYgBOk/dRmOR7JcZqlwGKZk4wvNz/Be26RjuJSw1tzz/amvDewkGqs8h4R9nLm67wbh2JD
ED7ESXW9R1lFiDwu30IlEOosAiPt7qIoahzHzUI5G/8j6cMgp5ObRzT/qfA0lFmCyVXzsEuEdfm6
AO02I9q3QVz4QPAh/C7wtwqzU77YDlvsflirafcQwrYFIpVBZpZMIo1WThYpGmB9xszWIaT11ji9
slNB7Qhg5YaU0c/HSBDhuUIJFbmgU0JNIW7Z5xTm1o5U2u1BBFn5TxWUmuw/Xe9FYH2OHMCobfRo
bXH1pEjM0dZGohaOsQZFw4E6WE34vx9fJ67e8PKAjrbB+d75rYromVLz0ibWrUnXFlJJdVZqoKer
LLMNkkvxo/XH0tZcVmCOL2MCikaePPnm97jVlL1CF1mACZJeRmbgUnW2n0KVZ11b7bqDQ7FviqZI
p6gVEBRNjWDERIInl0kYqGBn2IAo/vUbhschABMp94jONTIKIvZmDbfMf1UmCEgC8J8pKNMrhIHW
Vcs9E6dqxKsMlXBqx5ixoP1U5bC+ak3AYqvA+CGcNTLWtm55/F00b1LcBQU51RzX9RgSeHou4GD3
hk+MR9UlcfvugPCFCa4DOED6/UCh9NvDPt/xsYxFWrX7ic2irk98ADahJzYGGKrQGHCL7L8dWUX9
Q1XgQYT73G82gzIeBTYJd666SMfNeUrnn0/3wQmomCps+NlwkqilF7QEfGucfPdFuCOSF5sH+rf6
WMzZ+fTGBqxoWatK5WaaUFpTQH9nuvZTwSfGZsAXLaiLZZjBPCMGCAX0OYF1URd6BoJubtylcFqz
65To1XXqvJv17nLDEWY0ZJRrFefxdg99Ne35EDEWKsC3ukYdccaIorLS1okAzHcEyPeEDpD34JC7
PB6UkRtp4xswANfVBVwBz1rQDB7sUB5vm+VQpm0mWm2nAPDmXaWxNYXDFf3aYerInXlIMpDY1BlI
HDqZwIiAKZuSYqXHNarXPuuQCXRXDRsoJxje1oudwDu5wbYFEzSYYA==
`protect end_protected
