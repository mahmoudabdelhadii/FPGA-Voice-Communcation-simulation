��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����N~@#�k�0!����+��=L���0�ԴZ�2�Mc���ZO�����=�����վ�	"cqw��a��TS[��{=:�����K��-�մ�(��k��N�-� 偙O��QZ��~rL'�x[�i,mׇp���O�I43��4d�,�H�����SN��d���3���r��m���̨T�I;uj2Y� Er�*p�Q$Gm���p�V�`�2^���,hz�<p��l�Bxt�5��s��\yq���#�@W���f:m��T�	,*�񞭋����_��㧋l�	�\�:��uGd��PǷ��N�I��_����Tuv� ���us�(H�~�{2H�:Zor�Q	#%�3ˠ!��iS��95�,?�.���/�F�i{#���Tp5����Ҥ0{%���2vpn���X�����@l����3dc�ק�3	�Ed&3�ZN O���z��s�yxӡt��v*}ԫy nj#��lc��m戭k[��5)�A#�����8�!�]�Z�s�M���t��w�!��'ÒE�rv��Ϝ�c@<U��\tq+��&|�&X1)C�����r�A~��B�&�����s�:n{p��͠R�X⺂L^��R����c���f��J^?��ܣR�O 1�rV���:��T�4���AD����˩�F�w��)Dm�O�b,�a���1$��c��7t[i2>�ޔ0,S���󧇳Ϟ�ᒨ�-��}�!6��Jyv�醊�^_�(�H�(y^����o#����X��3-�k\8�M�T�"`R�DF6ȕ� �,5�;Ҭ C�k���1\������k�t־9�}���� ���QHF��"��t�9 ?��{E_�7��!����](�S��0�q��w�9��=�i]�1�GʦȪc�W�XC�|�$��}q�6����zf(����լml�dz������*�eLD�*�,�m�]ہ6����D�Gw� �g��' A���FX��\өܹ&�6�h�Ð�$�(+��埧��= Eza ��찠pr[�c&��nP��x�2�TK�M�V���3Y4vIR\������ɭ�1՟?4�_y�y+����ƄJMm����@����m�����c�t�����:ud�Q�����T4���QxBŎ��\o���t�*Z�$�*7<�t~eP/`lfhg��6��[nn��#<����n�D:� ����4��� :P�L��{c==�G6���x�b���_D�e4�/��|�i�h#뤾��vB��V6��s��G���h��>܌���W��8��۹>��%%��K@>���{rVP{�?S�zms��,n]E������L�dG���K!�J�,JlʱtW?�m�D��c�B<����2�ߌ�( �̕Yc>-WRw?C1?�,�����e�.�ީ�Lb��z��Y�$+R�GS�Q����:㈋N��<w���RPW�CHC�h����WG]u�z_qA[ƿJ�����������5�g��PL4Xt��
,2�/E�)Ļ_f���F��hQI������0T�Γ>i{�I���&e>P/�����<D���F�V����8�M�$�Ȃ�U#�l�{C�{�j+D2U���V��#lC��F���p��fxd���W�K���|B�twS�[jB��{�%�e�w����Ke�!b�`��p���mb} ��5��5,�An��5�`Y#�ܺD�]��(pYl9L�������¼���cN�(F�ҳ��[񔗘/@f�M����,��!�`M��� ̝y�"�oݪ�\v���R�x($�锺�	_�
��%�x]A�*=s��r#1�H@j�J�v~����L�EI��F��eAV���˲-�8KN\��a�[��g�m��xO��aV�*�P4���L�s��Ѿ	q�wL��{��
����,�"4!�HJ���!���	�e�X�c#-�᳞��H��
�)�_�?0�{*(��f]b��@|��ӂ�������3yez��Ʃ5Mǯ
�43���H�i~�m�.P����M�0�	lZ7�r���M�j{2	�F�R�rZ>��H.a�*"ݘ�y��}:�`�7T������v���=�WK~)s�nZ���:���$����%v(��EgI�A����䴂�D�|�w_�pF9�j��1S�z�J�a���I���	��:МZ���n3GV��^�O�@�5��c�AS�awj��R�eP�[�E
�F�mQ7�b(���ه��&��&I�p�9��t�Jч������& :~���J`I������7|U��U~�O�P��m���f �F2m��S
�a�(=�w��0Q�a���J��h(�~�ː�{�m�t�����ѓ�=��}s$/4�/��n��:i�]���G��_ɜ�˻�+�x){�� �v���i��di���4�W�1�ӹv))u�����.�J���j���̓:f�*__��3R�7D?�;�S.�vb}�`�̽��?�ie�2_I��n6�����.�:�R��� 覰�i�Ҙ�~5g,}Λ�wH�iII���TP�?��K�|��
`��1��/2�i������<�&W��%}D�jk����]a��Yr���r��Б�-"M�኿b]2��q�e批�~՚d�������W+�`��#�Ml�=�����%7$�"7�$G*�E����`/����B.�0������.������Ȁ�\�<�e]y�����5ġ~��;�Q��j����D�8BR��S��*�� ]�+���-�Ϗ�rH��� ��!k�.j�|R�r31����7�C�q$�!�с��H�*m좺l�u�%C����T�� V��s��d��]w��ݞ<\�?������
}X�A�Yģ��� ��^v^��A�\�B�gn��_��W���+r,*mx��"!���K���ݰz�a��e.��k��`IƐY:0�#�c���6���3�����v�Z�f�$�P����G�I�\�]�z��̸-��(���=��K��y�þ��K�1��#��s5�|-x�Y���<�}|�Nz���^�X�W	�Ӄ���S��1�o%���3������i>���Hq	\��]���Y��u���)��6�ŉj^z�dᘒ;��lx�h������4�u.�7����;��5J����Z1B\!ܙg��M�W��[��4Ē��R�x��Ƨƅd��=wV�St��~�7`�0�%�6����N������"A��?moK� �BL?�����]�(�pVd�NgS��~��޵��������*���qԡo�h$�r��W���t��"ށ�_���2��c{`�R����t�'n�??k ����T�<����N;��P��e(KĒ�>C�u���.��u��VQa@�8�q\�R`tښf�PP�v7p'g��E`H.��:�L��>W�a�fLo��8�g��k���l�0W����U�wg}�#r�'b�pXvY�f��H�N���%�G�:މ$�M A �����x:�g^:u�/���YT̢^%���1��:�^�#�M��g2*��/8�=V�>��N�",7�����A�MS�������v������n%�'�Ұ��կ�>�*ۚ�^[��wI�n�$��I���I/i���hC%�Tw�� �7�����ʆ�� �m�q|,��K���9�u�wz�/%;��f4�N�h�;��K��U45�ʂ�VU���-���D��Q*+ܸ.9&�ec��()��c��>/G@fz�ڂD�Uve��{���S��	�k������h�ȫ=w|�9O)�ܨ��j�\��_�m�R��vpn�0����?��3bY���c�E߼�6�QE$P��G��V�T5��\���x�yS��#KY