-- (C) 2001-2016 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
eItw2l5nrErDfdEJQRHwA984EQYf/ERnuehodyOaqP7AoiobLkMiFt2entR1c+lSEiEOQEJckmiZ
B0BP5LBKhGdTIlpnj83a9Rcqc6vbPceOhSntC975wkFCukKoU/15AVjWbX9TQ9qoLs7JBfvWH6YR
blfERIz8+jYSmJ8oDAXqd7w1CCgHbuT1lzj6PhKaigdU5SKIYUg1OhDy2wJdVFUdCNLgUALW/Z5u
rvA5inBqgn9DE2dWdWY5JyMRPsJmG2MZz0YDPfv8vDIMt5JOH9GDoh/FhBOvalmNMOOmNzrhRcJY
WWdgz8mODoguw83/YmLTtchiTyj7H+LJH9dJVw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 20480)
`protect data_block
Gpqge+jzuO1RV++9SzRMG4MI5G24KuhszguuIaSjAV8l2KFJoQHBCLRuKLxhDQijlpq4kq/zAbW9
YbANPGzbbIQPEx63KkyJ9ev33bQt2M5Vm+0+uJtwqkWh8daf/yO5ff7lf3f/LpoPP/7wl12ePERL
CiU0svbR7ec6V+PK9u6AN30Rnobc9v97JgixxAI9ahdcMdaWsapR8S0sn0FOoxsA2fB2NNGJmR9q
qRJelOLDyKnccz1LnOrdJpzRvY+g0PbGSxOQreRMpbzwWsn4hAJpbOWN5oL8dqe5xBPHBjB3O4RP
bc2DmRvb2iiquuofalsZfv1bgzKFFjxqglUY5z+/V89iJo4VFQu1XGSbDKUNQhfoXsteY7FIUPih
RTzjoLsjWSYhjxVkw+/wDPKOHoS2w/TW438kdw5fMgjEfGrDROsm3q1rlf2hTQ3PyXMewv05DAaq
qzsWOrDMiCYO3JhkcZcSYrQiBy7VAxq/7aQ6Ok+X3coqy+OhOut30thXG1Ga0KJNCgG8HkpIotB4
gvHCp29n6xH9d7K+fqVNHkj8MREYiqbDU45Wif0yU8qgZv8LybguPqvZ5sM7PNoYHqZO2gjaoxme
TUcSBRQIF+1exrEHKz4wXF0HhMRxhFjLNOAKe6XnFbF6KZj7T4wMC1z+CUDfiqhJXLCOFYBXa7s9
rLSOIRGVN8LCpEJD+1GUEbFK5Dz8rCnk67xqTtYxe6dUSkfSn4I9AmlXZqN7V5hZHDpNj7IVlpWU
Pao5t/n/ghaPN8rwbAvAJDhmpuWcUn9iDACpIfsSJRdbdPy3L1axzZktfQh5WjEea3c75Pqj5UU1
+trSGkTBX2haCcm9NjSBYLHqvp48sUaKJZWBDLz948/rw3dJblVevHkN/NaQKgwKToQl2KQG8+Lk
KagWz+p3iHksYP6nOsTzoiTKFLqV411NLkmrnJANBm331iOBzyTQZHgmHnxuiMMUT0pIoQqSkG5v
L3626/zHymrhjMKDjSH60WHIDuQ/RAh4uSd7Aii0ber20VSEkd7e3HvGIMTBjKDqb1dp61Sj5XWT
sj4OwQ1sW1nA4kQec2IR5TO0lzfC5Cc9qX0gf07FmAxHiDKJglY0w8/CzwrNzT4pENekHcDA0IOr
CHgalcCuzAVbqnuThMU3SMAVCkN9p+piIjuLoK/pow0h2LrjRNx7s8z/NLoYOFGdQFQfL5pJTNcw
b2gOn0SWXfvr7QxvHTmiTaUTiwSJlpdssvxY6FUH0w1e/KPnyN2clDIPCnS1MrOzNjGjoQGVRps9
zZM9ViltQhTgXNR43P7MY1IVK19SnACWgK+kQMOcRykHM7RptXPSpq/8CZSJ27dAfkYH3nSvE+mr
VRlRBT1075mTZSdR5VuRnGN+6kqVfPbGiC9x7c/ViHMXeN/RtqG4c+jNTZopXzIBSCWAEmlXpCGx
cVV+QzEAVPir1uERb9aljQmIqO5x80RdY5HZ2U+11sFyORYZACRJym0t4UXskFYK88ljiXXcbo9y
84oBkRlL+pVuWOd/BxHH9LqETStAzangVVccvOh0D/XRkQQo7qlZLf7+uaRBapn/qRJdkzjlyuUZ
5LBksZ2SR9yZJmKi0Pavy3V+KK9KmRJEYzdJ+N9AdAGuMF1Vx4u+y/Cip9b4Awb1kSs8q5lXGSVW
gPDK7iTXV8/UNmjrG+b+AUQQ2a4gMf6voy/sNVVM5WCx/QJwSKLuT2EJfUl/9rwA3FsyXidKcqAL
35uyLo2JBE6s1j5BD1WEhyLVMiB71TWV7SlBUhGsMOqIfT0riyoYVUyEF5rLOaFqaQFyUqktU1Pi
Ip3k43kG3VEJSzx/hUE0jLJ2AHHS99JnrkoDgvyGldmUKcWlNfKlp1CLu8m8lI6/IQv2vgI2jXDf
PA+/3AEOTk6X/8hOuAG64E9sLPsOWYd9xC+cYBlUcxdwjleAZIi2RrqqZu+lGleY6ywIbHQQQnMi
RKzfGsjpxbAUy3gioHAIQ97r9ZajQIcTaYKegfcVPVDi/e6Mk4LElH6kIRLk1lLOoJFEza9ScX/0
9F61tnNjFjKLk/PXeMXHLKUTIKUqjWlSQptpBHfmT6YYOuD1yKZw9IfvB7IZyX9Xlgkrdo5f6HA4
v7uQi5aYi/9p69nRpp0YbjUx0ZG50jRpx9S/8vaqJE/H1LoiQbqeTliNEbqopdGVxQBqRiyBwVJS
EQz/tl9PbDG15YAMQx9dAZ9EwSu47/d8a/neG3A4n21xr6E/SU5yNTtxPPteQJtqf2V3Aqqs/lxf
3dx19aO76lDygWkLPODWRjFGcFnaoUL7HETQl1rmdaDWUuDVuccKmwTAp2h2+mfF7J/nM3JaGK1q
OGcvrTSxrLtFKLU7tdrMn7wcavuOtJEjw+YQnxG5f/6v8tHaZVvg/e15wAQQS8FTwKca3XKrA+eW
m7QkzzYIqVD416ALLa9p1qVDdqwPGNrpdkaoejyMj7lDGDO9Vdz1c6rMZtcsOVF/BDGhQs7GzG1u
NRYxeVRB9vPdCt6vXzW0m9GpYtT96x78Q4m2Hg6Ud6d4JbIAUD2QIUG+Hnebtqkrn5dqnwJjY744
fP5tNmNGJeLpr5h38IPc0cuDGNWDd3oz/zC5HdwLDSxbBweJhyvi1Kv9dyQTDau9lqEr0vE2juxY
vxJc2LgXbOBLAvRWXW9qQBZFe4BGA+wa7HKiZbvbkqcwn7/uyNIxj0e9uPg2cJiymVLfIsUfEFBG
cFlea5Qsr35shqY3gECbu+GURHbs20fpd3Hhk0fki4vbrIXfnR46zN3uqQ6SnhjP8zAJmv2GueJJ
jl813yK39d+lHIhL6Qx5Cc8GzZe5VmN8cvB9kiBdbVHYBJA1INwXbqvH7smNfD6I2VpPHGCbtCTc
Nlbwfr4UpQRfoHEuhenRijZsUisiPy9+JVfPjY9ZYG49u/N87qLziBmQUMRuoOzQNPevX8RNLCjN
P1rSTew0oe14Oqw2Mro6KopTpX9j6wyYFljIpWE9FjiH2bqONRz5MYd8RXLCqDHdMd2vmcplCdw5
l0rX5CYZCipukmle7+elOA4Lzq4xO9K4NCjJrkxMmMDJq36pq1YHe2h4nGuAbO6YN4MxnBs1DyOV
j/2BKhz0wvzl04qhbQrOaefJWJMtu29fkAHq6pRPSekukqgHu50/fQbPr0CdIOrqvU6wXs8HdDzy
SvyIHdDyOyn5HW2ZN//7VRndWWzOKeEurnXPxxFXkP+j/BPn/YdLm6DtCXEL5NLvc5AdvxI/TvIJ
+3JSZOLFLTxBvOCD+pA2xiEb/0LRtQzCALOYMoBuSb2+gVJHmJTOuSWp4IA3MtRKc23zbNBo1Azt
gTFsvhcKRLcFQLBddmuOs2/uDU3bioh/OTZdIMxLY4lk9LGuhkKz53UMvQ2VXMfBpsxA18iJYHUY
724Lkt5mgDwQZAXqCOCKcHAAWHeKqGqQ4C1ZT/tt/piD6CcG+ASMdM1EHHpGqLf9vKfl5W37fNSb
18Z6oUCQZnxI3CN/7cNYHrhGP5rf4iKGpuB+zeFbCXeujw1uIX4AAt+gw2rHxHi+RJuzHdTDIv76
tuMdeYTU7gYfXx+71glRsVfk/rYGJOJJa8Di4gdqnc8QuxWPBAipEk1l9QkiE46qkGaPBDN+vZ8D
1quYxWUYdHFH05THQ7AuSp7aNxXY8ZperAnwFDAXJZe5u0HAI0bzWah2rzziaBtty7xfto89OaTX
UJpaaOeNOmi7219Ef42+b9+YFe+WLuwZBbpU9ZsC1zeSfcYsS/x4aE0XXXkiB3uDolPZEUzpHHN2
EGrpl7yWrx5yrGh4DOgAMLlM3T5LFSwetmZU4yb67lVJZb/8NuEYae8M501qPAYvA8rvWjvAMQRP
Z/kj1+Li5crK2AnnIAgACSVgAsYeO7oRDeRs2lFpvBSs7L1Pa1ricHRXWKJCBLS7YIu4RAsXUcL9
WWDHWr0ehUZPPDlFBlGprs1kMrFjqjindFRxRlqihooSk1UFV/Cqm7ePG8ijprKyPGXTgAu8KfDR
T9TrdBIJP4ynGtmoaSahI4bf1F+RkbXlqcV96H+gY1OpOLYK0T8fxfrZ7252Pw5PbFdSBlcuIlmF
WB0yghyWq/IYUAxz8jmyal7Vwf7cE4LDjiHGeDLYFsrmaFnhI4so/jXZitT8xzwIP9qPGV62skTo
Q0iqZnrWd6tX5R09OiuP+510+DZDtIQq2wdv8qRqw8hYtgV2s4MPksoI+oUXKt2vZ4WWUv1oO2+t
MyUwDyRqx8YhQ/Qxm0LNWeZtO138nc8SbLyxLkOVxiuZKbQ9C3Id0r5K0V110ZRbD8rKjjR0lLN8
IZRFaoqDjk1CuhgpkE1eodCRq1R4Z8iHN5wDv3i/8Bv4eJ2GX0NiIqsT17Ys0LChhahU/qH/FYBk
6lQ1LE5uIm+QiUGy8MHFgz/vYbEyJlkSs5gzV4w3GxiZEg0DBiSqSE36MbPqoCodq+o2M+TEkhLr
oCjrBYD7+faBl6EXfCqOxgFpthnE/cKiTGTWamttfP5iWoEMyDhUS8XziKm6lV2K4ttFX+z793pU
o74cJa5AcqQHjZDJmQD7fZ8b8Eu3Wc5CCUseDMlvNzqZRGRAc95XLqkuuhit9SOI/5Mep9H8c6oK
WdXFbYedWk8Ky0XQW5RGvbSh7FIuxtubtnq5WD4gqkzgUhYgzWtMtMLY6l+kxdEhQsypglahBZHY
+w1TkqRPMTK3mAFjZ5WbshxcCDuqmHhZC7+NK1m93xi+h9SstNOFJzEOLNPaw374TYJzFvYR9a+c
t2TQ0PgUJzxQNAEDljPs5hqmBlaFHvPkjF6il7GpcBljLtof22CEe65ZTVG5jehYZ6TXzNRg3nXo
t9zk/MbK8dNxcAjlVMz64sedLOSPuzvzFDjx5ihfSD4id9MP67Ig4btK3Vfrb9BaUS9WAOENBXjz
pL4ffyG1tZ2DDtUIC4/TYrHyPusrxyVs/ZbkGl1QW3Q6MzQT8MHhxbPFdnHcl7R//+jIHxFEvV8a
x2NWlR5lp0DcZPygWfEstgDJ4GpJ8GKide0rNu0f7AzfaiGFegodFgZttC2H98zAJub9WPrbq0+6
OiACbE7ZxytuazPlnkw58LrSEU7f5PtnJP8Kua3NwPzPDyKQVZ+bAJR3jRFg6RfbjFiXRg3nbsIz
oFkVScOMaY3hzDC6JCDqTE6zDOZfwBNm4KQkD5vNVYq9e4b6G9tVjGyFG6AT9og+GVtF7Whpz7Rs
PlgI7Tyfci/ghAShiQ8G1PRGWqyueqyNXinL4CSa4bV0OowKZRMKAJQD+VJvkR8QL8af6ew0cRqJ
BUthnjEsiDbteJVFBlCWzksC8jhqqZyx6bxuKbAokgE28VkbhKP9JGo8huTwlbjqTbtP8hl7eMky
r26wT99zILHM1BxkXRXcUCjh0vwLqbjuq02qu4XWP8KcYsVex0Gbc7MeT0KOOcy8PZSQ1HWrc06s
4PCUMqgqguUaA3Fi/smN2xYWs2oB7dbLD50V/Ir1AWxryLH+wN7tkhrWYZV4qspDTv2tY6Uz38oD
ooPNDeIP0Gk/SeQo4LCXCi3cavZltMBVfu/sJtduRcgzR3Jt/K/yO6p0FVA79xqNlNWL3ZQ2SP8/
fJAUw6g4X0BDmcqA84HX8zEUrgqJYXCVl1anjJDdWOUR1qKzOhPJnZ48xRunsY0Tb8OD/kyTaSPg
wcxIQqu7n+UZFjXRxlb1FFRzTjjpLKRiwql4pWD8fpNb0KfhtBljqILTVHYg4cpRkA+4cKnozIoE
xphcHmaNkGXR+imKs2yVqLASYif1ETzSqEAeF59/ssjc6dc2VQ4CA2UlNJ2Gs/KqeXXs5NGWzIS/
RKk1lwcOGq4Sha3ZxvrnW5+AlzVRF7ISnKmbY/+7YDWrHc1mCeamZhjUdjfrvQHd7R5cblTEvXQZ
Rhjqh5DmgdXSi0owxMmMFdNieREHoxapgc9MWDTqCVwJ2XRTwrGIDrM6+e5wD2/bcZFSiFMsiLZv
P3W311FIUV6A7Zxf4m8F/Dw5EalYYwbj2pKHMEq5Cxwwn8YOGwyMpKn5Z0guDKH/NJSGX6rXslum
6ABmnnuhn9f7W/XYlgtSMQ+HwXW1qtShxIm/Nggy3E4ivNO9Dka/lSPFuvX1tksHOcHIyRYiUJgG
7d29dwLyRwX47IhOnOzVaPucLahg0bsKFmA4rDY3zYIe191/49PhXnBCJ1uH20HYgqRe5EO99NME
B5YfkrAcCAHyFKmqMUl8XgN0aSgvbZGslaSBLDxZrLNJVnrvFCIw706L9c2Igpb5qqSGMQ7MxF2b
NgmMu84s4xBZ+xv1LcS3lWYNoYGnXl3Rm4u00ee0i857RUOUJuAnRYDnwV3PBbNwpjAJqhOiB2vR
ZgQN4ZpB0xe577koH4yXfK8VQ0c+njkdEUcmrPHt6AyGC2YKUBYP2OU6a0kxpJ0D6/WuXuu1rfHs
SI8AEXT4xpWjrlQXZL8h52XetSmiIFAhPrRdFLIv/M6jP36AkzDGqrIG+wwvsmHv+4+H0vUKIOhh
QeJb8k1cEDR26sCxIb51YQKj6cPw+QkuiTIoGNtaGPRNmeSd8+8jdnBel/hAwOmGjRm5yHo63U+9
MOs/Gnbr5mlZ726gi3LEzxSNdZXjf717Hkj1fZrMtjdXx+ehU3XDKtTPTeQO9mfiHzbCM/lH+sHo
CHcHzl7zBkbg0Z6edJ5h4xN95SaIXuVORVbaJUxoHnw9JONTIEbppIWYsArOPx1GoMSiquJ5wAyz
clRywHdOY65m6IDWLPPgECLQdV5e4YhifvXyZw3MQ/kp6vXxIzMHQxzK90v6P77icJ9ECFkXnopm
oVUccF240OKjD4tCWL6+JBRMJj1svmxDEMulc1DvlcMciW3QUGncL9V1YkSaUFbjslYgfSMomdx4
tC6kOMwvGEYeNrRE81sGj5e8xf6vbUHcXO+WyA4luDsgnuzm148+vSrqyIn43IeypCBE/FD30/l4
3Oa9nWLO2tFLRhXoPWDmWchj6SUhsCI9EC1hMUgdlbOe62Ql5+SDld+QTuqQT3MDsxfBO7wqiKCl
V5xdS0Ip007ks8HSkMilEJREI4MUVbVacGChzNIx47ScX8Ie/G7tU9LYlW7aSRYLWO7Lk8aaqN4W
TDzyWJ781KZRcRV7r56tBYReBktAkqPTdN1QfTvkriSD+ZaIzKt/Aol6dwWwm66Xpj2qlDZF97An
+iMrLuAmFD40iR5xTZc1lxpMml39p9Brlf+bUIRRr2Yh8tY/SW390q+fvWbNhXzRLAKBcMMhgDsF
KaE4hXl7KGXPtAjRBahtizSophgJj4Og3CDOhYeMxB7gBacK5zDFhSJ23kFBH137RfEUw5HV2sSE
4TraH8QfbPySkQ7RE5h1iAAfCmFANn3VwR1NvTM/KiTesL7tLM6ke+M+5bjPL01gYdJP0G1JEi19
cDkgeEE4fNpF2aqswhS8vXHWe5L4Dzs+p4KpxMHr6Mr2EuH45/YbIZCR3GDedi2YEPksyKqQ4aCH
Tx9djM5RIQ3hVcP7K9uDunYG2NhZaJfdpRuGekL62tiSWeC3tfOwWfLdcmhQiT1HnfBfva9UkjKt
1hnTOiZ699wnq3lwdAijRhRI7E6ckZa1k6cNynvYqibXPkFDUMjOGXctIOh8kE7aUjhbYgMfxdQm
HONv4n9UxoHtKxItLAiw1bjpBgzHwB7/lxfdcNIwNWdkPWnNm/htBEeJUVQtrRcLp3mjIi1nSXOk
RIH7M2nrtJP95NW/01Ua0timppXTgCN/i4Y9hhDImv6tbvrwb+mnlFhAe1jrTRaMRUMa0g/pSkaA
ZABi5Fql76wPTrDGj9/rj7YLpAa6vv+7dzdXSJoeQm7k+LCQRlzFct7vCQt11qxXitNJ22+nJ+WC
JqVm5kNUu/dZZZtYHEGh7HvXAhb4scKAH1QlEVmzY3SV0EvrDEX96jT5JUcMgg3NmDlcTLgcC72W
0m9kELofoex3f20LncBHsoDZHtmdwMM7+RqTdZhygudDFfG9GNS43yjPsXFxrI0qgSq0Vw/b2OXN
yXrdGzNzWJl1VXO+YZfC1jehJUocVqIcl2v+xUA796DPvM1dc4vUhEoiZApIgnZVBw5Fac8tTxfm
6QmKFK+InABr+IiVicByQyCOU4K2IECKj6VtvrdNxh57UfTOQhTURDHoMoaEgGIxfDcRusOlMsaF
2gc9Vi/jFFn6Ry8be2wpStqIgR1e195kRcT9AsJgAOqo5rEBH3KZ9JlU0bIYyFHCUh1eu53oqrrC
/Bs6/xJJ42ol01VYQlAUmHyZ0WarBBb08Cz8/sztfnpbuLBAXcvJYw414s6admjWv12iFWyycZle
f4+/u3SpGix35XngjSnEXjEF4k4Jn1pEXhOe8A4CAigbTh/fhxb4FrrvHN9XAwkhjpElNgeh39/W
/20FajhJMlb/ZD9T0zPKuU3CoDRv77GLx4whEU2LZatE0UPRwSRAglBGvTc4vmHP595353lKS+3h
3SMZon9FkdNmMN4NLO8XFYA0QEaDgE7V1guJCsu2rsaNwKjImQ4x4KNj522pTurl8AkbRhb/Xv4z
5cJj4RrwrslRNq3aIoiGn5z1iyoED2/eWwzGp6j2hd72h5yGE0Ax1xksvPX663x9imP4VQvzBTbp
tkWdo8m37Ow09iovD8yhlt93fNaxDITbKZEZEiY+i6q5Ic68POrtFPTDWqsSW5PLwYtxn6kH8Gui
U41bz2GOKRVERhUHRx6VkbGapgtNP+oi6u+/SfaSbj50w7VVV0wvrrZ7KFtJ9vOUJr+1aQQ7Z4eN
eIL4wZVhJOKd+DrR75ZMiOrcgaF3dM8Hs4M5B7AkBqQ3Avx1EOiuRMd04/v8lmyvvrjSgIH324IJ
l60sl9UJLVgHE+f+Cb4UgT8B0kgvMmqOod6hj3I7IEWGI4VSZY3b2vNntCQrec0e3UgrF/GEizWE
ctruFLIoiyqm3dBhThNqKTgq04vIBt5Uor9a0xoxwiuk5QrDgqYvc0V2MmzJ1CKyKZ4JSWN/bgs2
7UNLNMT0UB1jpvDEDuJnB6QTBHF6ZgQaoQcwrQtp06M1GY7m7Ez4/UWis9H6bYk5+7Y60ppy5Dco
nnoyoIM/wUF6uuLiYUnE+kfUAlXBdE8Mf3GKLjHUd19vx7ADnxtd5AV8Rly97DiYFk3x0qA7EjBc
gz1UxOVn7nsxWYG2y5dTvjYVhVpgnRyA7ayrYCZAhZQaP36AV9OuulFfL6fo9xdFNPLLLulZf3T7
fawKbAwrvaOpfX+oO6eghRUxcLAK8rYMGFdjONKx6fIL8CzkvGlHLnPQE2hfjWIeYMuuYCLqpL3l
7Bo+ecAzGGe7x4J8UM1rRTvcHYJGsXi7wxg5CeTiLu7NzFq6g+loQZj92K3cxBAx+eN4XPyWw2XK
EyhYsKNJXO8WZrCzJMWag4ChoL/rVXz279RGkSsud1lvHHZP+CxL9eapENawaIOMFEoyJYMDVWD7
vVDJZZPVRHFH+/SymgR7p5ayZxmlc5lVVSFiZIX+YjybNJu4GkE4eDGbTH0qDNVkbc1mL+FbtMvu
qIEAVrHSNIVojaLZBkrQBCY2+BOqX/Pm2ddS4/NZhRlTjhgh5K1sTumis/QUtrJJ2Hrfh4kWAQHT
NSx3qiPiEIddFc+2msqHDxyIKxQujmVgekw6maDHLgr3fHndwLpl7IRKz5uHOfGNkhmoGzu6HIIT
TLY/Axi9NilQdB2zL6jmw1Uq5yLjCGCghNPj/n+jwNeA2dQujpgpXSil9qGx0+gR/dXzwF47vMxx
x2uBAilPn02bBwxYWtXmm7frZeKhRA5v4vU0VK8qf7tFRU4aeyzAOiSL+HJfbrBQyJYGlcQSO6IF
6wuBPdu8tLpKOYFIq2FogZgxfzlQHSqU2ZPykGGaMHlf7z1QRuzMAFHG4c+Iwopp3PUlNHv956NC
vcOS8ifg8Yvx9J6D+oogyOk9Wu/UDxxkkDkNhx1IVpY+LC9EiDZx+Pf4ItMserg85wO2mmF88zWH
RhizcvPNBagKX+2hSdWGw+eQeRC1/I3IUBP0Psa4eCUEyEjDNXA6yh34MzS0JDbn+ssKHbKrv0DM
C2tD40Axbev5no4l0lM3zuoaSX4CVBnYpa2vyrmqtPoewNGU9BFJizX90kEDLNBIstBM0ePzCUtE
hYkl+PIcrqiIoWR8aPHriJdNC6/E3k0g1081r/JYzxxlKdWYAntmovfeePaCSjWVWHSJWtTZgEVF
HCCyFGY4YZ67lP8kmv3Z6lL809+eaU+6f0FuXI1KTSTrE/cs8jTdZPYSsUm0mAfLRuP+G7D3+umX
17R6TSE2JG2FptmLVXr0Gvk6Ydvrd2u75ZgyjJCKcE1MF9N5B0OD/+fOeopm0WYVo7wMzJE6gKA/
tqCyhobAQb0wPPmnNd49si3KDwJdBAwy5/uGYFGCOaNFhAh3ivdrw/X0GyTd7gwk3Le0QHe3tT3J
Ff8oREra30StB7DpYLAKGZcKYde3BacnB0uoU40qHqB2exj6HFsCAl8fZU5hdyyYJPog4U4SOJ9z
AFRbTbFQKGC8kzF/Kpsb9p2sztlZr1v9GXTG20y83RUpile9egenXhd5yOVoAa9olUOyTvB8I0Oy
6kIEndeOG0pcjaHd1Qbx0GOPe1rmAe5pwUgxeuVKuANqLnfg3jsEhYZMJIKyUrLQB6ahJNoZZDpp
Lu+7zCfApuGfVee2EbKVRraYtM9vw00oeP2R31GejaK8r84GIJC1LSKFhGu8kHrDdJL6v+Yp/xxR
iJ4M1687D6dS0XO8Mk/lai372jYkkaqVodIMnxGU6H4wI1U0DdcNlsacokdHTN4CxZkgp8VyJPgB
712Yws/uYPdlsLPcB6RFnwKfv74bH36AawncssD7rECjBSozLgZKZaIPbU8gt95ojd/vC/wnh72i
WG3EgeqXd80QsLkcJ8vk/igM3KDrZAQn7Y5THG8OyvQ8z2czm4D0hWuHaX7zOaH1e+F1XmbWe9E7
vJ/87e9VRVb0Jw7cnoPsLamCoFvH9zNCmkg0BRXRXyXH8qg24LzEiUWZ+3FKHRQdHVQLkb0Sbk+V
2iyHj7dfYRNfYO623JAaS4gAB6dLbmLLKWBDgCjhmBFB3+Zo/xrQmByD/RObPZ7V1hMU+/S3kE4B
KTvw8Jmyw1MWb+0iWGW93uQeVyZl6+B+igvZnuk20wqQK6XqNU87nGXhKj6gki0qmu5dHlEP7Jgp
s+7eUNRvsr1NRN2FUCprZ1Bvleiy3SxNkNko8CZ/8Bca7r0VMJr1mOQN6ifOjp4ceYN5BapaY9Np
/yE8eqRNuoMFz7HmT7qDOf6Oi6X/hzfsKCv1aO+/onjXxXuzR9NLNOsqPZ66A8cQvbn6mXVTLJ8t
5ms4JIKR7WImsqDCmXEIMpccckzYlIbQ3oYOgblIt6KDiH/aFseaL1tXJRJvwg0xA5dj9/Zm09Bl
T2rqr+hAtESYJ3NfM+wTCYrri6SjovgKk60yajuLl6OFIBH6vSJEY0W8Rj4Q+7hDSqSKh93VgZHu
RiaVIU8zjAGeboXlY/98s2nNQx0OO6wdKEu+EkhUtM8HnQwVB3+Hxu7vIf1GG4yMBpoTKMhUst0i
OI9LSE1ohTWnZwnyk+qwzrO6uqpjga/ZxEh9VgyFY1kMtyhzeUcetfUB9xqB2CDLZuZrtmOMlfpj
x2EXCqy2GS08uZwErAmGWj9uXKSwCKGnX26METgB8wsTwkuNx9UqtT7A+pzfPRxvUO4MmWZ03N4X
0c56SR2kMkYyFyyjse1+4XVs3bxYqxhVlugrbhjVM2jnhZYqUx5VEOo7bkLW4eOnzP8+6i1ku7SY
Ly0f2BTQD8He9RadhHIudbYWxE3qmBPhQPe63cdR/rcRx6G50jmhnu59MnqGvGkY0HzROltP4HOv
RwWQ8rFd8JJgfGuz3e96x0HEIwAUmGMzLhAm9tBha3x85Pu/qe5IFHnXVuAH1rtMm+enKMjRV26x
gBrTP0qkur7v/ofyJ6jPYdspGMG/WroLfTNajjvOVzA3mmZ8PQhbQQu0APNEKG5Ie7CsLcAx5MCa
lQ5GWWdfyLVN28SJKTPm1VpNdrq2iJygEQRjrp1sxSn5dUB4WQR1JH9rWTqCtKUZIljZHOPKlcuT
UgmzontUn8tqYFK77pr7I7XO99O9H18XfWv/IcgPAmf/QNS7Hq75C6CBBeCooSCLfU1rulshQXZu
9VeFcDSvpwL1rllbhcaLMR1BvfSjdo8Q+Y5ndp2Nyfz11qezLm2+xpOGxNKRoMIc9sgzsH+XNP0e
6sL8e8mfomDpapIFCE72I1o/SsHErnAHt3QwskwQuB4WuOLne6d0iakBotBB6NFN7OlG3CBJ49OO
VixhPjd+XbNq8uAIRdsmd3aZBRFRb0ErZsZq1GzXUNFMIx3uLWH5e/RcQdQSn5A1K22IXL2Em6TY
/PHqZhTqOHUaPlZ9CNGxToigtohFwAAf8HpTrKkHhuPHPrbELhN+VTmRmNGQK2sazMuR8/gBl9g+
SXdw6HevRWb+DC12SIoYXroxvFCq0Qt4dQVn2OmGDZUaOEZ0wvwKZj7wk3yrEgMthAeDWY85oklx
98CH7uP/gI2XGuB5Vq2oh4uGrKAePrFKEpt4qbs4ypqJm/nwvswerPzTDPJQTnRYdAdhGhjzG9Ft
7r3/rJYnqV6p8KrXOkGcu6k33bd5RibWbgCl6Ue+/pBBZ2o28Qok7bApTu5PWyn3PMP9dOICeUFT
rOWL+mvK3vtWsnaYApkXxe7NrhiaLMSiOgu/VL0ZEAa8T0Lb6CtciM3FgFzZQ90joP3EYh/IEv6z
RlrYRA0B7VGyZGa8v41wbWwcgGZIYuUgr5QB98CKnDReMIxZwkkwyUORW0oZa2IT6xooaOOciE7+
R0iDYTEbldJ5knkU+mvtCNQZA2vUhgckPiOA16ZGSgrSZyEB8QvAxiotytNTACtwNpRX1FHLjNeu
Er3iti76I/sdbD7vCn6oGTLgHWdXROmQK9tj+L4bdeBaBoLzCrxIcVmO0rUKjDK74BnygC45RILk
QlXhnbapI5QC1J+2vdBpw4xIZBrSTG7LRoo62iHE8Sd/AjTHOXfuqxIfiMDzT0zq4yxMsodV3u8/
2XuCVTV7tM3Hl6Emg/gdeGZlJ3w4iB2+UI1BPoOT8ytUHgoK//uSSONegH/rj+Z3zt8rhV01sVKP
eXIBjBMqVk/xuDYQUtMPqbgiVnFdeynP2GdEcu57SehbAg1ilw3/mLIKgt9NJNonZpycjJNIgqtE
LgrYyDMIy6+hg4zEp650LwqasbaUbNVXyiZpN7yD+/nmKW7u7HlDZ7r7Jy2Q3M8m2LabTtB+N4Vy
QqCWXnviz3pRKfSxHQJRjeNtNc7NWvI0Xj+n1rl2F6idqL6qiUMTOz3WRFPHbOLwRW7bS0aroG7Q
Ghqa2Rrii6+sPKiGANxp75BkxqBf9qzB1JCibHAVNGZcL3ygZB42tuoE2h+Fb1dJfanm9RREgwb1
DE92aWesi5U8GIpQFTU+hqnCSJ64s36L48lh2DtaPgCpoSUJGIdf3nbzohNhcK/1QSlngLHsVXTe
RDH4c7CMt5OjZUp+0Zffv/lVI6qLMOixMeWhK00PSmT93g9/pBEbC3UMH+zKVS3oQEn3d6BDmyWo
EAMSqLJaMuD/+CZtRwnwDI9XeHtYhb+guBCS/q8mZQ7issqX4Q+A1rskPUNsfnWtyhN7gpGp0R7c
rZ67j4czyF79sgPHqnUY/W77GhdVWTSUkcXZq8n5NA5DaCcVNt2RYUfKt/8DntxP4Bf919lGN/5m
RDGk1GvdDFfaenP+ej/aOEqmzPG0QKmH/cG64hfsA8u8jXhisIvOmqBwxdOjOuP2GxiKmJsgyiS9
Jlqj7tn5k1VUEBXsEIs77EbyJL/TY6xqKY4+SwH6JRE29y04/Q1Ysqpa64zATc7ue6EGsDl6SRjo
FoLT7Z0cTJ1Jg5mSbbBt60Y3TDeh7kh0Of8eVC7UaZcTkBs9EAgQ2BeFdYBN49R2FlSw2CQS89VE
f0g15XrdGoSkoLgxOm3awqhnLWZYEGbq2KUNly5k+8FnI/Em5s1eMEq3kM0nf4I0sDAaw81tAlf8
5PXF6PF8CYYaBV/alD9rXfc9q8ge9JBkQcE/DrLnrfuQcI42YAU6abHL/SkJneLPXMZE6mXF36bs
6liHIH3a1HkdT5vFAWHhW9IbXb4Httu0NuN8kBo9FGJFKezENppoak+3BIJZ1XPjOKs/XLCZw9QS
TAuItTaY+cEJOAEFZN8Z/4P+ZldSPaWFgBaU6vWQTpDFXCLdsUOQWBGYgOczI3ztcgGNnkvu757c
zQRDq+sBBppHrDyE1XwM/GfYLiEPnz8HJQDvzGAu+KUplV24VzFfGs6PR6Nn/SRwN8HgSKA5a/h0
gQ91zh73gD+74K2dOStiw7bqiSjxqFfT/YU9QE0A0VM0Ocs5KpBGpBoKaM9QCugq184VUI3X5ATj
xZEAXu1nYCLo4Vs8MkIX4jmGXHVp0+w3kaeJuLqpcyT22+Uf2wK9jxci4W6mOBkf/SnqgkaLljQu
mLalouFERtOqTgtstImIjlC2zc3QhleYfbX84JWL2FrXlIDp3sL9J65vQQFfN+Ciom9gUr4s9aZW
K8ptQdUG8HL/ZV0lzrLycc0VV1tUdHc6eM/8gVjIbGajCwB7Lrf1I2tVyt4qdul66g+NMjZfZ8SD
BrW/ZSD36wpbeOHNSgZyfKYOFgbbdPmGaOlVZ5XVh0ROhDILLi1pF+euLLSURDDbjYSQqRBB1/G4
tLLx8cZB3ur3QvKEa2NK5j7+mlDjeuG+tquqOwbzn0siIT+nHKguDf+O3EQqGkNbfl8rSGH/vQqA
OUD22WzBQdi8GXgMu3aXQ62PdirXeu57VuSCMvbvILz4JxlZBNwxMmKEzM8HXcNwxs6fi7o6sO8k
TcMZX8gt9fQV3qAvZ7Ab3rPdyx46+zKDWLRxbe8xY7C72rfJpLJzoZjOg3ieiFfDEAlRedb/0+tL
qJDG38zrCrc2gZpO8oAyv1xRWhcsDeKGtM0mBCJ6l0nKlGrwwJA1lTWBEjDDztSVLGJ9LgQEXl90
n8gjQ0IvoL/E4plJO60PAqbfHykBOcuvYMGP9rhih+XbUVDGsdPteY/KPCD4Gij8eN4/RarthxJY
qbmYCVlnQhtADOhn/T8NnAAYnfJG42v3t2J7Q4Pfm7OoDVPWMamANG9FFvQUgkmwnaQMCa4S8A+c
0SZO2M5MxL3xaX6moV9TiWnZ3F9OiEkMSNwNK6fw/O3U/a145dWfRMiQQtppDqjqfXxFUUjLqKFJ
JfNIQrHFX+1ai7JMA5fY+1LmxwzuT0caVO6B2pxUYrV324No4V+/F/+hFhkwi3GKCFxqbZ++6U1d
Vq/vslz2Le1BefL8bYfFVn1RQlEvtjPksEEMqSZLcl0Vocc8+DcTfS80pErd7tS+yurbPc8NHCBx
9oYmmszcirxFJ8TwI2TNgH6nShyRlvHGv+HNDtyYTAdQ15xizjx8m73LElEH7zuuzEl4KDKeyyUw
4uRg8OJ/gJOYJbkUqN2uEGHmATJE6f3zj6DF7jZu4y++Ge1oXhBka3WUexFOdhmUMYXKb28OC5gr
Y4tnkDAsI2XGKeSUgAYKN4xtL/uX0jSYPdcP9aEi17EtdDyXhhgzgzR4rBiZX1rvX2BgKB1i5i+0
CFjSWc2eYR0OhPW8X2XD2KLhP4cWf/Ze9YEwYvAb5ogfxoP5p7ANTZpc6timhilwXHEvz00Lu4Of
TudXgoVfIZYBfeGnbvjFVicoq8Ga70+PMuEtKXo7JfcRTVngeBDCcxgwf0nfy3STnksQ6kmtDQGJ
PSy932BzgNJaIYOu+zrfYv1H9SF/m7iyqQYpI6PPgV6mSesLE89eIEc/cHzS5Ygq8CNi84SGR4Pa
jGQV6h6+JSfgWo7Zk+lgCPN6yaxmxYEWgxkaWv9azXRD3vNsxkEd9GbcSdK4YyqeT16HpI81DLi3
a/fD9hFAMBk5zk23SVfDEFr/IoPTDMqO8CZd/onHJwFm7XRQ8KQg0r6O8/cRCzkt12RpW0toUMlO
FnOoJ33sUwRXR1TSVZ304cYvizEvpar2IgY5Fw29P635O3yPPv4WU8uP8Xbm78B8w+I92IeRL/Cu
vxPFWy9gc6n71HvQsNKV/YQVoVOM5lCBLAy5a6yOK9aGfQvyiliObxp3nf/kmPRPL0ArwjLfYQ8U
vFRk387Nc1pNsfcraF/zmLvE7tsC7i81rDBENHsc9+BhBr3n0QlhXbz12A9xoSUILm6q68BBrph9
CSEYlTrasqbbKzwTagxYOaI/Ng9TqYitk3mrVuwmoFV8uL3JgfdU0Mngssg7DUDOFjczAGQ3rVyY
a/6bv4ygWf2cYTmj36+eyic9bEpJ4BxT8bVg2KysqiGiwQcWlU0ydxUvtTLKUp6dP+J9ndT7lltV
1CiDK6lDdJhuEMq7YoH1T6l5xmRkYgLC7X6C/KoYe+YG5M/RWbY1+M4cTUMFluTefmrY13XGyglY
HTUh/cCtYnl7BTDJHWM8xPi5ygtCrOfN47zugoid+xEpwdkEy+HoLGQJa5a7/IIpoyLPvEqWGBSF
UwLyjnBZyEmHinHs4T57qUad1VQ/JlfknqWtJfEk7J0Kmpt6mwgkRPwxIChhilsZfgU1PK5u+u3e
rcqP/Mt1HAOJer5ERhoKstt2UynXf11UM7QodOoWK4CRsUW295nAlo5XYuPjwFdEOw29fhsa4kcU
HjjUlF6gLYFbOoCwn14JRHttrM6xAqAVH4ejAEnaHZp950YGH2FTS+/PBzvtOokwC0afMKYdmbMP
S6npLfk/p1guCJ0AL3GIjd+aCIpf2kCpGGup9Jt9wEALJsZrIiJhwgvinfKFkDdBxMe3XcxFS036
FXMtX9bnmyZ1IHN032MSYIMRn/WINDyneGtzemt2dpOcHEk78IQjlM7IGboNMV7TjFJNEMHg9Tp4
uK9wBklyuhfIRiN8cEPMi8GvsXcilZx9Jz84wbLgmQwCu4GqcgYuo87wI58n+b96jeDnKqj5uGEI
8FEcK/L/NBPhT3K5qDYcegeJ2ZUtez5HyD+wJby6HqmrDsXKEjj6rnLKtL/uV5UfwnNZs6v9t5h6
z/73f+vhsUj+ADFNzqg7xOfXFLC2UVa2JUEwXdDJYT2z5zhUfzEMKb+03UqvvoQ6Gzj+et83iw/5
xiFJHrANxd0/k88KkfTKeNxv94OEZvb5zuT1DaJsW9bCHtKss43c1+ooGvBQMTktf+IctLQCqEbg
sKWLMp3dIPnXeUOSCZ9UlNv1jt5q42l2FQNcNoLWtO9yK96YLC+mnxCPheRy5WfBbFBMnhafhRzz
rUB8kJEtFLiF/WeugdX9Z5e02iOEcvWCGEFTGtp+2ZcDVvdL7U4xmZTSH5eX/bIV9UxOkUV4cQVh
nQH/5d8V1pYy/m3NQPZSBfnarYHvAEl/fsxz6eygxDsLftM5CJT0qelKDcmRaBHrtbzPZflmZKGF
4JoNg1lKhZSlBAoemqbOEGJ+iV6EpgUdHw3liGpQSqgdOZZaYRoslkIsQa+5Nxe8uI/hvru+4zfs
d1bHrjPBYd0zfH3aE3ZWIC9YVsLUKqd/wX2jiMMd0peSTnY9zoZTZvShl0H9eM0amPpyQlkqGPpw
z1sz6Hl81jonkkwjhQ7noqwyRVks6zk8ImrRfOKqEAIipSgJ3Hyc3b/nflxOtyWLshltV3HePU//
IO6m3fv5KPDaSpehVaUr1TTfcSFjAuBeI+pZZA5Z16wCBqP6OrQiaQTRhBAvE+Qt+lylCMZFfF5G
G9Wg8Oa1VrMMRNJN711ciKrSIuvioGvhap0b28mvPmHh/fGkMc1BkW7yWjX30tyN5r4d1f5F9ubC
0pcVXX+t/4jX+Q2Qxr1bqmZ1Q4XpIzQLl4sDRCGVxyBWDZ/5iaD01tlfSU5rfPGOxW7xAKrpIDFE
ZN5q9c2GMQlakINVAxUmaRV2UcQULus/EXjHzDZyY35Uf0zaZH+lu66xa03PIPtt8ZFJoNnFYqk2
y2etlbJ3GjGiPHIvI+ynMeBLjNQsZS23/UBrUW0TEz/SjTvRMVyDYApuFxc2i2FMBaEvCVyJrkJT
vHSljPx6qlCuW3toWx0n470JLtEXtbb23B0BAjciGm/ubDxtXOFNHsCG/AgCDeZjALyap8zsuybP
ZzMeLOImBxhBIvruBrfUs+VoXDDivfaVOfcA93U8s9jE1C0VUNejLtIXc7j3O2BFtvs2tJrelx7l
t9AZq8MaHwfKcqFWH8TrcyTW0XP7HlZ86X6d3ILZKomdUxHtRt9U0+MSGUpKQfx4H96VfeA66uQ8
xdehh7woijUqkzs9HnlvJAoIjcX+jT2YJ4BWzyxbrCFI2iTt0yV2b/lapKuaIe2S6+qGsq73p23f
QA8bm0MM1j3qLA5os319ugExtBZlx8r9EvurdScsXrNYMV3jVlBjTb3TORxuC1XT0DYatuGGDCre
6VZ5vFUpWL03xXOt5vjkqPIn3g4wXJy2rWkaWwMnernV5bTzvLmdivSl3LIhWhN0ksODAOpCExju
vwUiTXs0HhoUku4IziuRtc14CbkXLpF7Rg4E+ajOyhiJHC5IdEDW6UROZhaHtfagFC1AkF83CD2D
/EUpWwRrmE6LAN4c7KsIRtEDm3nZF0APpHkacgcI3zPE8sQvkqM+Y8BxvMoNI6DWT+fIqvgmcToO
0gnL1jObt9aJSpUE6k+78oBu3ruShAjkDJNM32lP2a3b15eoSN+SAwG5x5dmfkTdNFMcMJcxFi6u
IbDdY6BX5Tt7hvBNAtiH6UydhU0osjHrNtxQ12ApnmadsEFnPo1VXLKLBxtxPfGoY6yy/oL7yPCz
/JpuBBXEN1p9KayGdMMkNgWWW0P55aBrOz6bU6o/JepAI09NTRdxZii3/zUrXmwI+Wymy7cS6WO1
+hZ5jUV/ggGbU602OhElE96pNGh11eRQndKQCUjwtan+BdXLOjBulcqkeafnlODiel6HDom/qb91
8Md6KN4Z0E9ZXr2SGDcoX0YmtDrLpBnREGI42GH2T8vtbwUwIljHmNNL/wJj7wNkiKDQq/7o4GG1
a47dfZKY/PIXA2/4zrY/NwY676ayz4gtxQGfJaMv8Jd455f406QCls0G8BPNThI7QMXOydPDr6Wh
oS+e9qnXPyjmzotOc6DNUPKOW5g+pGUEPgHNazRER9yqjvxNCxUR62vNPStsknuhQMRPazJYGZIz
vGMsoQemjGlG5hJgUl3XRbGa1BL4Jc4oSv4TX14GYL2SP7LVYFYE2xsVQibNgNOSPtYs6qWp6Z3e
FjTD8wmnX9bCYJ+0ZBbkqmdgjg0M7EpOGelPBcJwKKLblGRWwbBs0lrhH8GtbnlGivkqIZ8B3P+m
aDlS9oMp486NGJj8ee+aoLxhU53gQoHd2TOZZGHdgCz5KnrL+mX0BYs137w8fLk+UBsg/kah15NL
2fYCZYOWiqDr3Al4OOIjXhbHHY9xTYfJZPinaLKA6FXsLU0GAYtrrLTDMZDKwULmoP595ikWe7P8
1Jz+aOSbXAIMTT87znUbFj1NuN9bNMnNoakUQuS93HaMbEgA5RIzHI5Nc3yp4UZbjED00UIUe3yA
HMbXfFAflxIzQL4RKLoa7k4pbiLsCaxvIm4FrSd4QSkYoVY0ybnOVXi8ZfEdaAqn5hNZlOqSI8xL
fupkc+OZ28oRfZpaXAE5yqQVgR2BsosBtW2UH+FJKIqZ5AokiaOrtBVBcGqpW77kMj4VZw22RtL/
aw7gE332iJXwNT4I90YzCVu/hvzdMu6lk8/snIeER2IxP4z7asX9xfW9MeC23EdqYOh2mLTmTyED
md0SBAznQ7WP0ma5gYA3P4WhPcYkAjXoYDouHYpCs+XRKUF5h626WoVYRIMVT2lK70h5PQ7Ekmm5
F1e+zKb1XrzVAykNLboFWiJJtRNQlOybbP/7anvekRJ4VsYgKGdo/KmjHnxz1WRF1Nlenyh6LEO2
POQrsCqMCTtmhSHUPNvx9SOWKX3bO52wwDOK1e5mjN+W22BPIFB1XeEo7uPRpYWTeq+J5XnzDKx0
1DRk2Q5cL5P06SYMgWNTZnfCeS+dYT4mSpFDWVEXl/I+wnnrCrUJjkqCH/2V5v7qwD0tDptaGXZl
afWzzVj9Y64YLd7lSBx497vTEKkIQ7DQklZJ8TmiNYcFnRLvQH/GOxMf85NcRKr0g5REdfH8NvGo
Twnivt6DS+Anar14mItzBDeLeSYsZRC6p/BAlEbU/f2BgZ1w8e7Yfn7zw55GpQnNV5BL+c0ZXuzS
IeNioMeeaUPfC8JbVt7/qZil0JpAy6qU34drUV688FkqoniKY/y5pV1oGzkGgh1jnXxI0qdEs3ws
AygTr0OPn+sb1mBvX07UOLvWghpas4ci5yuLE6wtG6XFJHrDKVe5+sSc6q4V5pt/jyQ716ZtetzC
QvEimT+fO5pf25ihpwsz6H6AgZUbavXKy6U5WQhed2z+TqgNWKyuhSR5f+skIRn7qUVoA72QZYht
cVvHTJk1YtylM8SjEUGY8mEBr+pUC5OxX8hPAjEsP9AMa7j/pKQ+tJb2ILB7Duh2hP3YAD7ob1B/
PYQTjDJPUuHSAizzXDoIYFudyvnC8EV1kRzPIG66kTd8Qm144xyjTTKTV4ATXqqbzCuhuJgD3EnM
1EPw8WzU2Ou2KZ6XOnIs/RVbRsfyZqSWf5S2Qftil3HumKxvTuDOzbgg5nbdiq8wlMM+gJ54L4is
zW6nilXVu6LyR1hIHK9SF6VKtsW3tHUWIOFINbhN4pTyMlCDow5R7bsnrm1geNSfIwRMqIXwIs4B
oQ82ypV/idD4dbq4MMVd58EbWJcTpmH+rD6HYupXBSC9UlcASCufXePBRBvwefiM96x3jcgdoCA1
yOMt94VrwC/Pa4hHWG0vodyYqKf87j2AZDvpsa/chSnnKGWvAEeC0q08uRwU+7PjIuHBBA/sRi1k
U3aOsh0eGzOJ0TipojgQ3cq0YahPP0NMCKwPxHhGJg7427/Br3/3TMQXc9F6GCJAb9jvBS1xS0XI
qE1wjg5DSdqvpHpasYug5qPkf0LNC5O08W0gehV6y79p2pUYJfGAn7POkqvXR4IdkaZGwNBlruZw
Ttv+n50O4hqU8yTzJGJDuXjWjTiQXfZ4jBpjsjsxrRA3ggi5lpyUj5LDIc1LRNvz74vE5uWLSjFr
BJmtRtLEFrtidWmy4DHrwZluaXxGaDEUksTo6CTy0YS2z63Kn3ZZ1UnM1nirAiKzttIRpc3kW0Vx
S7RI2/EG36UuMHfLF8/q9QL+elVEoQn/4LKCQ8DO/MI5kZf2JHbytvaCcRC94SEqH9p3FKOe0ze+
LQj4fre+Jw3q84iPF8AQ1eVC/h9Yzxr0rt7RlhDW8xP88/yV078aDK0Vz32Gvvhfi0kN9JDVFOJu
9Nsu/ZO4pYY/CnDt3x9728yVLJdESD0baiORWV1jNflBB3m6f5M0QSuG52s5SFjLXyaJo7a4yxGB
67AUlD31s/naQhq128xBXFvP3Gf3mt+77s33VuuYgE/KprOoSdiAyB+X6jPcBDb1lPQ8MT+s8+IA
qo6nJCqv+EAigUCfF72Bjs9YobeGEEZTMQBchzJvoEjZtQ8YQd17+MW1JZChvwX1Vn42xOBHCO8K
TXiQS5MsQEAqjWHn01k4bm+wPEaf2i0AUW8Z7cWWm8km8gAc/pRR4jb7Bz6eSzH6Xf8B5nmtOX8C
ORAV1latlye0VCkvIaL5UKrbo3DYgWvUV0ywdXnHoFH1XIJGQLPoa5BILAhHPcQHp9oOQC8B5Bly
QAaPTAjhrw3D5pQM3hRkUFWY4vHOMIwxuZir0C3TukP/MRBvAXcfUvpcdS76JAZLRGWTR242eeOJ
oBywH77evxTAqA5hdYkvAyVbcBMmSXshSOt81mnnnFcVHJotjAcCFE7zhyjJ9e2n/tmanLPo17b2
QdsU86flT13VfUAuj8I9+z9vn19q52WPdilP1EVswpJ6KFOFY87GT6TytJ0aQVihXWXKEup9AveI
OAjE7SJe6zNVvMIHQTBBmvxTGPn9hXdzGRvLcfkA7QRy2Bh5r4y8U0VkFo/qjHqgo1t/CzjQGfJ+
BB313hKyOUCLhh9BumPx3d+vCR3XVRQlSV7HgKeNR4y0R5fXa6rjlm5fyiWABHG79c6mY2iLIeLy
VGm9vOKl5BJMppr1zl7dYYzZfAUIvtM1Tde4TTdF75KyfAcnNjynR/3+0S+Qimmwuy6foTq+oPcA
TWsYH2cUm0qfXmap9lFpqTA7593Dn+vYl4EO9w+cgW7GfJKT9eLkMeo8q03IRYM7mbQKte/RZ4xe
SXF1T3LCBhxZv7gKV6RY56uM2Ia2JG72llUYtMQXNV1GS+nhC6Wau18PdIf0I09Jdd+EiE2bu6yJ
phGYlQU90UiN67W6F6zwxbBDtRreTC563VPCcM31/sV6HgRmdd86TbKVRTQNI9jKi0dwh1kDwwpC
PEFcwS5sUtX2U4Fv8BK7JEiEQQUZ6L/16ITDBwh8bslF2QWH7SVvSBDpKM+/1K22GIxJTs8Tvx9p
c2N/O/kCvG4Qv9cVPzh+I1WPgv/dMIcoBsLiP0Km0S8+MQI4JC3fTvmQHlsTl/w8vp0zLIC3i5l1
v8HfaT3PUHtJ7a9otu1Fxqi7BNXRJo8EGrplAYj9Cf7mMO8fk3v0qCBXDhtxqSZUkbQIZOh3xGeu
0OIUhnssKs8Mm6tKU+R/bfP75/iUQ1f8gibsILypInOZaYvlLQYbbNp1cD0uCRjtjrfG3hwK1G5F
hn4pa5slx+VCIpUVA7CPGPAiaobBADUFW7maKhR1AUzy6jCleXswOPdUSAO5THQVu5Hn2LIc0L8i
b293UVLeKOs5zKoJ3hCScMA1hm7MnUmdDygymtYO4bsFRIrzaKH8O0doDi5BOTqpwMuVyZT7NOIa
UqVkWZvwpnuVOvSexDC+sr2MxEE7xSfBaYKIr9OAqKGpsCuScwi1ZvmMz69o4X+hgY0Tj2x+sbq1
wKm9E1krNBZn9eosnsAGN0HmYfJaFEWW/lQsqxuCshCr/QXA7PzC0SDOc43TTlA0XNT9R+zSnvP/
Mz+hP+ouLVBt04NhGKHEtM++vmUzPWUZ46x4+hjWalJrIPX0K9vtvIJogEdhtwkeoSU5Em/Uej+j
n1vvVhOExnw3PZPCkWittlLljrkxK+2TjCUM/LQOC92OQv1ZUHZgQxoB3Z0tgJwBkKaeGVknX/AQ
Q0nsyJd15YvgudST882CMt6++l0CYEn6WXHD+K3YcLBr7Eat04+san6m7fY/gmuGfzVag1ojL8va
ZgZsNTR4XRwe17i9GwiJNuml7Ucv6VYTqaACaUBInjF6doDFaV1d5nGrnyZqSitHGcwfttWBLaYQ
MoelCuLuZL2+k5wsnKQ+jv22oqB+BxP0FAn5+bhfGvx8Ppdx2Olg4Z4jvxMfVWoP1XkM1DET2Ybn
ECIMuI9yLFq1kVLbk0lfT41wqSe6mVPOFDOBGMnAYJv1tI6n20SD5eZELmMJTu5G/tOwCsvHgbkT
QUcEuPuKZ3ebLDsQGatCYwC4fVAOgq+CtpTvAlzlvLj7DZOmJht+MU/OVQF9topJDScA0npjoRMX
rZwlW9AuiZNFcWdvr5wrC1oYazQObCTSMP34xkNkhLAy/2uugR10vU9wQw+u8+P2E8f1+QnctMw4
uQRDcpjlIE2xxRHr0rIKhs0csJrMaH6jUgwJO7Fb0XICqx00EeU2dW5JYSB2bW2lGWknTnIkU4B1
xp0PGwse5jqp6itMwYKrnVeB5+Svp1TmmgPeJxroejRzg/I9aewvnM/mjhcTLt3AHjlP7KtEzm6z
5j8MnC1uPpQmFpbrI7lS/izWIYabhxXZ6qStHzH6MKqkgf25wL5EzAGCU+5GWHt0sjefhDvqMNSl
JK+x08r7NTYzxzbEDy5cy9vka0tnvpdy66u1uZNQg5h+roiS9rETP2H1dUFv0EPOXJplpIcUWWcL
TF5FQ4bGe3V7FFPJ3TBuhNGt6+BHh397JALFK0w1SV42zmsamk4tSAVSwEGHunYQie2yXera9w6b
jIR/0HTY2g8j8HThyFm+XUjEAdPD1AyTs7EfS7t2ydlxNin0jI0Oc9S9P6pnTB9z5GrqNf9Ie7Fq
RMmOUk4Vvv19PjplJ71hJMBofhfO/hml0uB8fY21t70nUtNPp+taczsylSXtiqBZAvE1VmxMNU9i
ZP7ZUsC5hmKZkgoQHiK2tQiEUE9BoxrxvJrE89rCi/aX5i3axozU2m6L5rzd72t9l34l59OxhSjh
LWMv1kTnVy2wOLPUNClr9PLhZr8wlA2vKu8vyrrP8wq9APUjYTqBjxkl219W29hsgQFl21mV9BDX
2KRNDAa13504umDs6iHCcDC5ei622gNqwhVajzCq3z9ba0jHz3nybWgdoUMmf/ctyOip7OjwaScE
ltls54XkRCgrAMAa1id/GwzvCm+05IPfOK2v4Zyc0OYYJl8cSGTsrfN/bNX2aDOOsC4M2E7Sva2X
MJRkpbqMqFiuIbaV7I9/EIZgAnbtdYGOnHQLqeiXssh82dk6KVZDczdKwIB4chjKlCfACBzYA6Kx
lYSGhe0YpI1O1jAJNLPuloSr4129fA+r7nFwTMJuBhvyanjg6ObMUmUC21QiP9efxKH3vjD1TKRf
i+p2OJwCd10ZuyK1cHfE0u6LeQFY+9hx7c/WBBaFu7iVIGyBkaditDZNaI6Ste2CnSM/g+G2xI4d
e9nTEXLgRCpW8UgaIgbkFTXAtWrBHlGs0X8lOyJDaYLb7z32rGiy9MG8yZm2/kqcv718NGRdLjze
yHjU5SrEIwPWGmC2id24tjZtVLqHdbu6iyaOX/Xh4ehZT5mUU+5pDuTAkpO0+g6SGHhZr0mPxvRv
8/D+1ALzr9rX2+KZ39vl3rpCvp1ywqv1mcyhF8AMzOZnaWSV2ruxCPjlZbl1K1uiyLoufnEn4i/8
y2MhtUkhCckCPGfhjCa30LWGQPB/Evyz9lInSvdvITYdtlNVyG9WWc06I1WVD7KphAtsvPkvUqIK
gOwj7co4CIzWxafl0JHvsZNZceSbUfbvJdNVW0vK2RueqUPy8+9hCmFUmrkHciSlxQiPtbDLCXPS
pDaI5dbnbGRJI21Y1JdDFRtLsLkcOesgbJ/ZaAUJsTBbX4V6FKSNrxAGJgKNY+YpVoN5+0fsEB5+
VztMcShuHqiauyMZiVwur8P7LCZDh1oQDuBKYioYKIf/9y2S4HFzAzdG4G0E7SigkqQ21558X+q3
aYcOBYLcut0x3jzIUg5vWmHFHyskZEWk4SFGxcKMov1tF8FmWcG0syRbwxU3cdfGTQeEJOLO2Jzr
gvfmZsm5PHte093aCke9Te0IjeyGiGFD5R2dpDzkBt28Ta7p82begAQy1KMXTVW16I3VNIK/NuOz
39x7ktC9Y9p/OZgdHYLZ7Z4rqpl8BukxIKzcGSKtFEANNA2JYrrFomnnKGH8LAjqg1GdRV/klSyA
x8M3SOuJkbY45YMMRj+Fn7d93jzhGlwkJeMr9X0U4Y5OBrFXkucD6EeFWCKle076Et4ytJGfUxda
unE4YHl4k7N6DQS3ro/6dcgl+DoqKlbHwbFhLY4r8hkrzWdglWTVqiJRIstmT+N3qzh8vG1qo6Px
T9EZNMlcrMDQMr6LUgFiNlLrxEwkftTJ+zCSyV5pQto4HCDk+xuc4SfLBf2rJjGctoMVhLeWFgwQ
phUoyjc5BVlNgM7mvXCEC6wcfUrWbXCzdNSoMxS2FO/Hea3+aMAux8d89uoFNNLirnRwUV2JmDEv
L46XmGRuoToW4LkdmbXh62yGTb1v0va4NivqGHiSt2t+Fy1Mx3MKXyf1BgyVdmSBnmvrrvJELsjs
zdhKqWRT5CDOx4mQ2fo2ovUyXQvaXAi6aSqfvUhfbZQByrgixEJVG8aDNvKW+rLhyvhJ8cxBLAUH
qN6vCurIpCB2yBNzb3aNxUOFKz6VJNfgrdkjw5KinWb0TsK9XhNWIjaiL34A/Kuynd31rNfag0Q2
PIalub7DioU+azx2dlDMNVTBX6jVv2PMgOf0E2tVwkolKL9aDI5D1nbq5qjOH27cxuI1vFtyOOaI
Ts4qUCzF2tD+mtegDksFDfurWXZFp0VvKOI3y3gH06Ddf8VWzSP8ZWMukU+JUPSx2mWwqjDOrF4E
9wr8yXTk8hWnXj1GqLHTvwk/xLHuAMHUaKwvYC1a2hcj2sLc8RKY2DFEFeC8aUrbVwmwIP7F8dC8
+MD6FQuI7dz7unH+wwuRTWskkvd3NchuEYhCcCMgDn0WkmubLr1arkPXL/gBmlc+X9KWjYggdZmo
Iseh5sS1F7QAL9TBq/vf1rmZclMegrjuJTGbgaaHyVchRaSc4Am1UXfecomF/DPEx+LpVg9O8FMS
n9fNSawX22QeS6+4idlapdVwTooEcw2lC2qlRCybrtTuciJ1OjHA3x/v2TGqgB17Ouuhyp5Va0hI
43q8x6cKx7A/OCl8ELWX+ckYAlkRigd0ilZ6zldLnSm8+aF8rNzYI8GD0Jc2iuDhbbStexfOrmR7
/fDys1SS3SVZv/k8WUCO4x8eQTqslF6OvTU0Cba9jUJwmiiG2LNPNwCg77PfjRQvVrshHhQdIEsL
1PqkgpwxYE8vn9KiAA8s1TwUSiTskGxpM8LqfbCOiT4n1OPMxjbP2aDwsfSkPjZ97eZ1oyBJ97JR
55PZi9GXYxjtkBmAzHiizhAhWqvqvGFGwkYdspqPOjdrONyAu2ELNTvSCB7kgOXFgmQkFLWPjLlD
VvxM5VObzMDLJ7daInCkzne1/0U9nx96LuT0DCk94/cjfLy9T8d0LlhAuNjVXBeuLZaTVh2lvQll
UmRQkL/yMx/o0eQl7shMik1yj38dtHZ6VAXDQI3kIwGVco00jtq+d9jejceuxvG8z1bGpWPKvWAC
yFy3Zsm7OX9sV/ezA92cdvDYdNqGYcUO4jZWzcoYqqyLjAwsJKM6NQXKzI2Cy4dSsoNPqG3Y9vdN
WV0uSnbEPkzDbvCvKzmuYzVD0zqbt4m4yGUWsykmhUslqA348K8l1NS7AzLGKGYg4WNklSkZNUQe
p9QbDHWjAhCYMHcRa5N+L0lhoc2f9FbDaC6Wy1IoUMJs+1+j0rSx+AiLMjXeNA7ScRyA4OkUAPLy
Ir50HCSGFS1uNsQ9oeNBxoE=
`protect end_protected
