��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��,�y�}�ǰ�=4d�H���`I"��W�`r���T:tB�T4D�m�)�	1��I�t��
��8(�8t>s)ו�."[�漆���]�~�]��;�O(1#5�-� 偙O��QZ��~rL'�x[�i,mׇp���O�I43��4d�,�H�����SN��d���3���r��m���̨T�I;uj2Y� Er�*p�Q$Gm���p�V�`�2^���,hz�<p��l�Bxt�5��s��\yq���#�@W���f:m��T�	,*�񞭋����_��㧋l�	�\�:��uGd��PǷ��N�I��_����Tuv� ���us�(H�~�{2H�:Zor�Q	#%�3ˠ!��iS��95�,?�.���/�F�i{#���Tp5����Ҥ0{%���2vpn���X�����@l����3dc�ק�3	�Ed&3�ZN O���z��s�yxӡt��v*}ԫy nj#��lc��m戭k[��5)�A#�����8�!�]�Z�s�M���t��w�!��'ÒE�rv��Ϝ�c@<U��\tq+��&|�&X1)C�����r�A~��B�&�����s�:n{p��͠R�X⺂L^��R����c���f��J^?��ܣR�O 1�rV���:��T�4���AD����˩�F�w��)Dm�O�b,�a���1$��c��7t[i2>�ޔ0,S���󧇳Ϟ�ᒨ�-��}�!6��Jyv�醊�^_�(�H�(y^����o#����X��3-�k\8�M�T�"`R�DF6ȕ� �,5�;Ҭ C�k���1\������k�t־9�}���� ���QHF��"��t�9 ?��{E_�7��!����](�S��0�q��w�9��=�i]�1�GʦȪc�W�XC�|�$��}q�6����zf(����լml�dz������*�eLD�*�,�m�]ہ6����D�Gw� �g��' A��)�m���b��ӎ���o�6ūvO��=�W�������}��	����z
��z�&�P�K#�^Qץ�_������&�)�ٺ�u#uD�	' �/|�qf�M&P)�tL�x�?�u�����ҽ�����*c"q/�\��YDl2n֢�vtX��Q������ǰ�6K�gVL��ο��Q�������-�˚e��"gb�_� L01�D��ثU�8-��Nw�@�$[�>V,���6�����=����{>G6��v�����φ+Y��	�d�A��b<�)��Gp���k�(�vWu����!5Y�N�z<V�<���".�����2L��s���`������6�<�U�Q���I,�l��@�xH)�����v�_B����~����J���񚣶�;_w8z��?g��v���%H?\]d	۩q��¦�6xIo#�λ`6Jy�����;E�(o)咫������4���h�� H�nU�5��6�?Z�+�jݼ2�����-��+#�g	TAS�
���� ]��_�6ڨ�^�b�[=*��7�fQ��z�&a��ظw����s�k~�;+��K`�K6D��-��#�UJA��f��a��t�����L���G����@?��*�|��%+J�h1�ɾP�'��m���_T�>�;+�.���Ya���E��CR�^{��-l'L���ԡ�N�{bR�d9g{�~ ��e�rI[;Ǳ֬"��W����E�-��²����4�2��~.g���c�yjc�-���}�
r���H�U�����;���^0��R*�O��N
�Äc�N�{����WU�׍�:��&��@Hԅ��g��T5���s��>1���:�7�L�R����,]�C�	�d#R�?ǩ�L�� qvC�"�τ���$��R��Hw\�|2���S ��L�Yz$�ؐ�E}f���@y�&�����p�B�6��m�7�s�S[��H�6��7��~�s��I�|	��������|�xL�?����~_#�*+��9��Ϝ\�{$�,#�u�ʗ�4T@�����wJ3������6�GZ*!����Ng��"6t:p,sʾ`�?��
E/��UV���ٖ��g@��"ΝM�o�տSL:�3��d�jY�AS5� �r���@ ��J��[Jm�ހ��6o�sd��`oåC`���5K�U�r&�+e���F �n`=ivM,n$K7�K~���IO����Q拗��rc}v��-��~���� �rبM�r��o.S�����n��r���Uә4tK�!i���waJ�%p��k�qs�ga�@y���@`&J�?���~�%�e|��xW\�In:vp����ג>6���p-w*�5ھ�>�֕	[�$������.�����.ltp�PĎ�N��S�Y)
y�^�ޞ�V@�Aw�Ԗ �zEQ����@�h�"���[�̖p׹���0Wn>��r��?ԥ��; k��_���=�q�,��#�#�w��Pz�0���фtd�2E��֎{T�7�2A�72���j���t(�o�)=�Pu5�3��Hx?��x�y���@�?���;��/�+�jxB��$wK��jWJ����[���������'�8����R|� �X����N�R�7$��g��R"e��-�A�_�䑞<����F�l��7��z.��߃�֫hۨ���Q؉Z��)k�u;�ɦ��[�Ƌ��ig��dN�t��!��'�)ձ��������r��P�]��<�)����������2pK7P��TI��И�tb��Lm���|�-�w��"�%���krQ�^����)M��_�{E���]�. YK�kB���ŖƊ�/�m&\�3��^![v�̉�cO+����{�Yp�<����� ��6)bƒıPQJ�ɻ �"���k�cJz���[+cs���O_0�"����������q��]]�oF�<m
:4�I�JԚu�fP�슀�]MrV�z�g�h��1o.f�ޱ�Fo	{<8ǰ���i���U�u�"�/\�;����S�0���Q�N@B�%yz���}U_�u|n��9�³�!l�jφ=k6`}<o�zA���m!�!㸗���}����ɝ5PȌ8�] .�k�p�#�2�;�H���7e(�4�D��r�,Y�2'��+4�#r�mi
&yE���G����(���p���1�vY���Xc�����s��@3�������;�-L��k�>1��Q�2�N��q��}��#ذ��l}V�WǓ�v��\�}"WZx���'D�!�Lp�4W��aI�7���Mqb�v��^��5*�B�<n����ഢ�iu��4������62��@����J�S��S�Ј���}�ӜqF��V{&�I� �ש�C68j���{U��K]Bƶ{�&ׅ-;�>K����"҉)"��t��!��UKąZ^�b�o��h,���.
N#���sИ�O����
>���"�rQ�������F�Ġ�BY����5Cby4u.���Z�`K��OY���.��d������O�̑�L�0�d�ºkGe��#I�i9TO$D`�l�5
�M�a(���+f<w��4N��9%���]��1�4�j���� �?
�nR��E��X,���~���n,�ֶ�����rG!h�8/�����,����
!K 7p��^�%�pf�<c[c�!p��z4��#�����ߧ����������7<��#Uӑ$�{tB����T�[B�J'���2N��O逿p��Ϧ�2Y�iJ���i�[u��U����`��r���^��3w�L�ox4A&��+�s��uY�*�Y�w��L���f�2�fTEv���_�4�/��ρ�z"H�i�ϖp�8}ؓ�R
1p�n% ++�lp�H�=W�M�H�����Ɗqd;�D�t��
�C�4ۏ��rhAv�Ps�v|�%��}��Ա�r�K�2}E���
-Ӎ�~o(��S	�(t`.��H�"N�vB#[��A��Z���&��~�$_�ݬ�+-���F��(ʶj>��}����"\�e��������l��JA}k)t����Ќ����1p0���6���\�	��&��4=�+��N'8�ঠ��<��/���ʇ8��	I���/��G`�ŗ?L3x|�
Uψ«jR�'v�F��-t^i��ߊ5�$y���0v��o!�]�}�w�3��$�<�=$Pz�2i�"Bb��&��`�ܶw�d ��a������%/G��w���G"tG�_�~����Ձm���5nB9�	aH��9O��pK]X�����*��S�[�GFMT��Z�n52��lƖ�hQ*ڹ����	���Z��±^'̋o�[�?d��^:��I�*��� ��|*���+%���v����|�/�Ӎ?�*��[E6����V5���`6�iXY��$�yYZ���HP���eNЃ���p$FP�!4�Nirk�]��8�+uDeF<-1n'X�E8�:p�c���XG�����IL��ˇ�J�nׂ��+2�ҝ��T:�+D~� ��I��hq[4J�Oɱ��23�".�E˚���Tg���ہ�0�U��G`5�D�s������)Y�e(W
��M�D���#|}�s���/����Ɠczk��,���}"�IN7����#�<<s\�]M>�RC'o���`4������ј
�@I�)M�ba��%A��sR����n@׾����eT�&h�H����1������ŹI��Q+
d��q���rL�տn��Z���_����D�E�%5A��Gr�nP������NZD�i�����t�X��8�>%8�ţ���eo�O}R���W`�;\*:06��oJ����s@����S�f7N߸���Қ}�b{�#N���Ͽ�������D��g���jp�if��c�-T-v%��I�Syܔ}2��2���E,_Gfc�>��e�c@(���@�2t/T꽇�s��<�h1�mM)�I��S|�Uצ���2�y�@�t�Ks���f����]@� ���%�uX�@Z�1un�ŃNk�?n�����O�!�����3���j�}�6w���%=E`�T!DP�Ƈ�d��5�~���i���N Mo�Q�u�����D�	 �	sV.k��8�!g"~�X�t�X�q�:w�Y�`��R頌@W��]/ڔI�M��[^�D������'����6�q��{-�8�Nc'|�8�DT�1��5�����]W|���$]f���g��ruB������d�\pᵂ��K!�U;i��k�ɓ��1P��&,�ο8���u/��� �"���g]������ �W��U)'��WSyl'[_�I�d���y��C2�A�_�	�N�lr��G�S	��[��z6@�yHا��7���q�l�����U�l |j�"K�~1�qXP?�BO$/�]�ݠ._��J��UhN�*��4�>���	�}S�Ai�,8�U�*h?sx`����%�Ω$p�bA�z�<O��(�j��	�bsX	�b�*�:z���|����J�(�l�B����~4��]'��`�����8>��w9V���V=�INb��d�^����<zv�f|�|=@��]
��+ؤJ ��v� ,��g��9=	���7Q�2R�r"����0�Zb���ۧH���xw���և��FP�����,�o�a��f�o�A�r�]*:�CDݒU�}��)�7���u���<+� 0��;�P5Ɩm��vk�t|g^�r7��h��y���PBϵ8\C����˟�_q�����v1i#�����W^Y��&_�v�f{�1�~93;ydo�2i7�\6`�M�Q���ƍ�I��Tt,��L�U�R\y�y�����.V�~�ڵ��<RO4D�ܭ8�u>�!|�!��!c���<��Z���,��;�"��u�qA��
�VԱ��~29�m��Y<�[� ��,�[N��&��7����jH����*@ܠ;�~�1����?�adv_Jre�b�-p&����硅+��6���)6�\��g�*hCd�C��H�u�Ro�f@���(�"��?�:���ԝ���6��Z޼����Im�с}�իJW��1�P`�L���/��#�~�<�c_��_�/.4���6���i��o�?㉤V�M�+y0��w�b��Ke�J��G�ɍ�DXa��?gq��n�{2n:g��{	/Ϛ��+}xe�H�sr2�wہϾ���ln{Q$�<G�!ind�FXs]U���Ң�@�����@#Ð�JW�*��hHJ�I����$����I��0��O�x��l^�E���0E����!,�E��Ѡ�V�d榩X_�m^\����e��紧�]
��\�LV00�_�]nZz#�z�,�o���.'`�Y��|��:4��ï�:d�yYǐ\�i6��A+�q�_�BA�H�U��V{�6|�oJ<�>?��`��:G=&}�Գ��S��LB��;�J5[��!Tx2S�%3H�93`Odi ��]y���9���W�ph�� <�vc��-!�U��Z~H�QYSvo���(���'D����n1;�BJ"����I�ռh��U�\�m�K.U33�ŉRn%Q�%�ń���ᘥ�F�Of���&�9h�v�!�/���%�PH-��h�V h �(�@�6/g2�:Y(�-G�3�~��)٪�%����ʒ�O�Y�+�J5��H/��q3�23J�%oF�q�_��JAԏ2�~n�6�6+�[6��#*�"��3�����\{�u.�-NVd�0y�t �i(���B���?=�C�
���:��$�J��$��C������"��g�C�4㭣����wK-�ac|�
~I��`Htú� ����6E����^���hQ�n��#��O//q�2��9���v�&�R�'���Ob �ns�����(��F��G*#�g���mdc��:)�x������ �0�P[��R�|�y,gh·��E�j��[T�ɴ������3R=;ǂ=������旱q�2ц�Z�~�w��T��68�7����E�Hf3I�o?��O��Bℋ�&WL��u��~ՙ��	YLڮʕ�������%$>��������d�i���~BêXZ�%�db���8�c���5�ޙ��)�8X*�K�>;�<�=��2��e��IZ��`ѓ�Z����Y����<~
÷�g�1B���c_�����XFn�F�K|�h[ G�mO1�"��WIt �[Ag�A�=_A�����@ �޽��]y������xt"K�%�F�e�Y�!Y���86T�յc�k�� �KvAV:��F����I����i2	^[u]g���] fÿ�B�ם�A�����m�D�&����pG��÷�7_?G�eha�)�T>��ɘ#O��"�Y��[x���t78ݑV�za��8�
ݦB�q�A'@���ڏ���!M��0D}�H愓�ܽ��~%�����k���;�b��M�VE�F���78XP{s:�pz�mW��̏��5���Ly�0�@
��)�������g	v�&��[0%����D�ƞR�r?ys��^�"���T�*��(~M��T!����"���o�NlV��r45���8������ajVeɢ���� �XI�sN}���F�<k�������E죽� ��46O�A�(�؅>�/d��*P�����N�)lk00����dH{>¸�]�!s4Q.g�t�e#���u���p;��%X�����ݥ���}*���(���Ho�^����"�]�1ߨ2!������6a��*����Y����uU���X�/s.�Ý�D�����6E�A��ͫ��ɍ �����t��lV�t�Zw�G��0OV�α%�W9�����#�^f�u~h�9��=��UT���+ EF������J�T��T&ALQ+t��k.Dzf��KжK	3�b���{��, �"��B���
�."�ˢ��;�H�D�}.�ȠE ��K��;z���.��qr�� �~�"�����w�����)B�٫�EM
�_��D,���?���)�8�-�
�u�fR���hG��
�i��>|�^�o�SY�k��_e.�|�FA(1�y�)��m<�@�د"�wy�GH������]�v#��dK"��<_� �x\v��J��;[�+��R���^�����
�N�����A�ј���d�@	k����U��#<s���a�I�w	��e�(z@�K����Y5�TCm|0HZ�r�e�D���l�sӠ[�fJ�96�#G|�)y�,����_+E����q�5pD ��e+�5Υ%D>�ֱɀ���;�汾���4�&�1���,��2���q�'�a,�TƗ��O�(�:��*�`�ܕ�����G|5?�r'�m�;JW�#?�[՘��X���ɾ �9\�D�W"~�{��,��p�7D��*�����D�����5D��Sn�O������H�HY�n�����i��yC7N�}-3�����h	����g�, ���&}( ����;�n!���ω��r���F�]�%(U�nr*�q�;���r�ne5���a>̷b��l+�u�t�Ȯ>���fw7$|)���M�&n�&Cq�(�8b|�y���EL�1sx}ѵ}�H�;��Y;������^�=�l$�RZ4ܥ�Eۡ��_�[���I�m����p�܌j�sQ�u1�vt^<a�K�F^�X,#��2�ڊ6���87=>�ǂ���`��8��<;tV7剗�~֗��Ž���R���톯`�����+�����N�L'���m ���� SȄ�ӧ�A��`Vp��wQ���!��,D���ݳ�.$�ʁߝ����5�^o�>�u^�l�3U��~-�Z;[���n0KD�P�����qfQHV�qUg`�{�Q==�=� �ڰ�Ǿ.*�!���0�Z����I5���s���,��&ֈG�W�5�e�<��WQ5�Z��nD��(��nɄ/+�I��4�=|0��MZ����d�&.<�+IA-�|�hp��U	�)���C.(Mn.A��j�({bo�I��0�XN�����Ǒ#��S95F�H���ׇ���m���j��w��g������u�6:��wk̕@��(#5��|�������H}�ԥ��̖2���d��W�'
B�YD�%?B�q8�J0��X�:�\ζ�s�C؉������p5`G�D��}װ�uY?zW@湶�D���R��E�N�ȱ��궨�I��Ժ�<<1?�,UR9o5�}�������|g�
堷����_�}��C2(h�*rۄ#�nu�)s�1|����=l�Η����s-�A���ǩ�ig���?��h���m�)�s��?;�Ē�%Q����;��f�a�� �������@���_�v��)n �u�&�2
z[�ri�BO��)T�ynFr��p������@P��h�������AN���i��8��C ��rE�o]U(����v�ؑ��W�h�)�'y#E%}��l�����5اD+���p=��(��j�avhl�z�T�Ky-Z^��V�6��W�
i=$�*}+_Eǟ�F�g���m��ݿ5��IA �>��ZW��Sl��Xu�0�s�%�34X�c�V�����᜞�IC��y�&e�>�B��̺�P
�L�V���>p��k�m�%�����)�3�kT?�N�y�OA`�G�.J�̡��퐹���w�����C�L��Iy��m�QY�#s��\�U��t凥��R�㓷~�cT�Ѹ
B�ѻi�L��Jv�����WOe��"�߄���-Y��A���+͆8w�r�@T�R�oU<k%�����N;�\��؂0�K{�z= ���ƫ�j���d0�̖�k�	&R}��4f0�S{�QcV%@-}5�9p�;X����� ��0NP:��-jwo����h�f>/$!I
��(k���0�~�q�S���Ә��q3VI�:����ނ/�'F�:���B��<L
������4��j)���Ӷ�G�('e[B߼+A~9ͤ�+e&5Q�H����%�6|$89�}����KW���dO��] ���'A�ٶ����l��$��$G^
��9C�2��zJ[_��Q�N}�b'�X@�"诚s[���5۽&E��՚��)��0�UK��b����"aS�)J<��ƒ�r�ᮿ�^��
�[@m�o��bi(T:��ju�^��v_��K�U�W̦׾�B���8���Lm!���/�����RaR���u?��2k���D�|CJ���`� �����ت�O�%�����<���FR�1��5kG�������5��@m�ŝF��m��6��O1UfC���%���@ϸ������%�p���9��x��Tf�B~ځ�Ww4T��$/o�?ZoEl/�$ ?�w�uZ��-Ry�~��j@o$^���Uc�ԡ��'�0����H%�h+�Y?3,��}���Z�؎� ���o�֚	�s@����;��D| >�c���@�G�C���P�H��ĵk��zB���>��ЛHZ�<{*��C!*7Qݸn�/�
2���I(�]���P}+�7�@����e��ď���A6��f�v��U2�ޑǟ���5wE��!4�N�K�'�(����fKY
��^I�9ki Z�۝�I��))��0��n3�U�䞗�2��LiG��	o�r�ħe+��|��vNnv	�i$�d���6���o9ј5geb�x`;b�q�8I�=%!�{L�-?3��ʄ�-�"��������h>�����
z4J�i��(Ehl�qg;�+L�Yɗk�5|�֊����r�`���ST��d�m��;N�d�UvfI�C=�,���lK�Ԉ{=Y��S$�����u�1�O��eS�5hD�^	���y��A挲W�Z]�y1�UC�'*�T��ߔش���d$;�mJ�ޖ����
?uwv�[-�Ac�q6���S �k����v~j����+_c�G���"���ׁ-�Z{�Z�n��\�H���q��\]���ޣi`P������h�b�Vpߞ�W����sR)�5�1��,�r���m����8]����FC|�D���y��;��@�Le�s-BW�
;o�،=�,F�f���&ⵃ��$	_L�ڑT��5���*t��_�� �(�S��8����{����Ǎ��հ��ܩ�]�]4��6l���U�Fު�ѵu�-/}d�ը����vV�!n�y����ɀR�O���Bdۓpl��-�Ts��-�]� AP�)<�7z@��>����RvQB,�����	��e%-&�5@�yv��o)q0��h�E�H������B�.n%&/K^�G�ʁO�ͅ�]i}��S���hLn�,���pi�b�u[�ٮL� ^�n����s�|ύt��Eȗ{k�A���� ��ө�.����S�M�p�� ���~�|�AN�)%���$����~j�4i��2��⚖,:/�����~bol������)]�>�j719�[���HՌ�����"�iP��R�W�6�U�X��m$�GNRGE��N&D� �#OV8��{�;��4;��޸���^�+��N�e5D϶/��IQ�!4��,����9��~jr1>��ofQ����pWX���t��f{�/&��A�xJ�!$p�]�O(�=����h�����T�H@Kq�D�M����-9�`����eL�g~r�q��Jwm� �ۇ��ݸ7�Km	�S�S�]�h�u�"#��9w�y?,ήhPja ��#/���6Rmg��&���F�����\�ެ��M�<�=�~�g
f�j8E�r0���Cs�Hˤ�6�)����S\��ؕ/o�t~�0#�9ޒ�r������<���?�7���s��!��)�F�q	ğ\�NV�I��D�����'C	�;�I{O53���똘:i�o1�4����X���1$8cBY �W��@36��^^1��0�8Yz`���k�.r�  �j����7y�)b&�.窃|GNwD���l#����Lnx\���`�aNE�D�X��<����]
�Z�uq��A�g���`�ܱ�,�엳b����\X�6�
���|���/�0�o+�4r�W��H+L�t��E��7�s���Uէd��CP8���5,?G?S�7s/2S���oB1���B����x��'~��l}�������22�IXW����	4��!�ӱ�hb�)�vx�t�/sO���7.���^i�?�:ϼ��v�m��kqI�p���$�b�'ơ����g*ՙ���pXQ8�K vк��~�����nk�P��9�i�A��%�rD����ŀ�+�e�V���b��3�b�`ĘL����,�X{d�+Ȼ^�O�@(�U�u��D�j'�Z�L@A`��48�A�7���snQ�;�.����v�;�@�YmL���0�u�����vm��UD��u]�/	l0��b��n�����h-V&�f/�3<��Z��5�&eN<h�ˢ�g�+��A����[�>E��� ��C��䥒��`,�AJ��ʎ=uZEFY��cI7�,9�{Yt�&�d􉐯�؆�x���3#�8���3Yf�n�c,*�%88S�"n��Z�~�a��4�z7�w|��~>j��U�6ɩ���4��z.1��K��v�L�۹�NzmJq�X+���E�&Q_�{ezS��`�g`��j>�	�9���@�u����s�JB�y�Y�Z�	Y���k�'��uI�#����J� s%� ���2 T�/1�M���G�ӂ\�S�Y2�n�6"�Y<\X���d�^���MIڎ=g~&a�wз:�_���x��i�Q�:���������p[����`�LoW�>�/�4����hI�@�\�����[V{�ƍ�~�
YP�G�1�=�Z��
�����.`�����Ng��}���N�Y��
����]IG���l���cm������qM+��|h>�46�c�N��R%F�t2#s��N�\o���9=��`��<l�������Q1��Kjb7��i��Z:Vw�UW܂[�<��3�Z�&"��_�l37ɗ�qO�G��ݾ��Z�	���>��	�4~Y�Z���kX5��\/�����w�,��$=��>���:����Hk��vd���EI5�u~
j�� ��]��N�&���`�(i�2��o�m��*�4MY[�J+������0�J��ꋝ$�!���}:�Z������4w�2�?(����"�i?� �&*/�Gr��Y�l^F������ac|NM�d�%�4��"���~$c2������T�}��Q��f3���ƤW8ܧ8nH5����������մ���[k�c�NI �+�hR�/�q]S��H��1=���n9zŉ��V�!y�n��n��E�� n�;�*�N�U���A�,�&����V>������V�Z̑r�iH��-N��@�,pY�.d���Q�>��� *��P,��4g}1Fz�Β�|VK�'{ۆB, �{��$�����w�ߓ->�����U2g3��o�K�7�&���x�(5=���ˀL�g��R��ʂ86|�n_�����͝hu}:��K]Go�Cxė�K�J�
2j�3�{0-�
�o����������_�P(3������f�����G����#7�;x���~b�C6�h������$)ꎭ,<�G����L�a)CZ\]�s�l�������%""@Y�p.��9pL��N�U��y$V�s	��=/ѫ�P��ל!<��σ���K'c E$�.�F����Eg�C��礰���}�r���
|���W�ȳ�l�.9���Ko���� z�S�Z��4�i���G�lg�k-N������Q������!]�ק!x&7�./��|�A�Z"�Rh�	!��-��[�O�$nl�$�!$v-Dd{�
�<���ބ�c���oC�U���O���u��2:�Qoi`0�������_!@�A8�b&�������^�6!Q�и��w�� ���3dV���Y&|XD����|���w��;ؿn��&�+�m')��?����*�Z�'�rQ~F�lQ� �4�	�J5���ΐy�$!L��q���ec\�����E���d.I����Q�*`�^��i�؞�gK�]�M��~{8R��O����J��3;�z��;��!48�QZ}n�xg����,ϫ�ʌ�bb���.:�C�q��5Ơ��˜��OGDY���W#m�ٰu,!A�n�p�go�~Q���%f�\��߮�2S�p����vZ�GY��X���{U��2�*�B��3�a
j��X�CL%lV��!ܤFg��?C��^:>��@j0Z(�hl@���X�.���բ���ͨ:���ϕW�ҙ��~��g �߈.9}+i��Uh
wLy���{�3�;� `��!Y�z�O笨����˿0C�Ÿ��'��@��;qrC�C����i�]��i�z��]h��^�z�Z��av?�h	����J<_0�}ӼV��!���k���q9���3�T��h��@�QK[=���Cٴ��vS0KtO�;hL�W{ҘE����rmOʣ�W��{�{�ށa��`�V?/th���$������5R�@<�$����Uv���O�����������68k5ho.��Jv�g��YZ.�jУ�#�X�ۍ�4^�B����g��= Z��(q���xZ',F]���Sj��:b�j�����(���R_��\�q�;�JÂ%Yڅ��� �&�3H���D0�G�u�8�ץA�k��˕���gug�E9!�]Ϟ��+���*���VYc.}�3Y6K�i�ao�0&��Pf�$	�0DB��D�TD-��p'��&C�99Q��3  n��u�y �4�I�㘏�|Z
��`ʶ�o$����@�|hke[�0|���]���%�f���'R��͇�(�0���L5�pfM�C"���	i{uP����S�	�P-�v	O�H=%n���.;1��Y���0���ߧt��W�~0��ʦj��î����iT,��50�3;���a8Yt>̐�87>ѭj?L���w�a���b�-J�E�F�hA���Ͽ�ngKGUr�n��f!.o����ƍ�O��`�Lm�~b��b�L��]׷��̙r(�{�,k\Urm�� /�˥��
�M�qs���zEc��A�ȵ�J������z������cp��T%jb�d��I�d������?ߚ�X�I����x��őI�{%��ЖGX�YC���W5+�ާ��v�܇�j�%y�<P��������i�$�%%�o�Ӏ����/,���z�x%1F���m�����.�щܵ�߼��`n�|�Fg9Q�a㴓>Y&�j����� ���"U�
{� qi�G�#>�<�~<U�g��b{It���(b	̖���ݯڋp��Vr���/�RK�j� �����y,�ŉ6;�N�@�Z��ПK���d�����9�]b���C�ٖ�t�L�)�R��c�����A3�>f�.�r�"����U�N��qa��8/�Sds�bp���cz��� �Q}?�$�a=��2�A�m���<���c�o�%��,>��fƲ1zo%Y���)rϥD���a6��\��j����Y_����xm�n>G�eL�b����wc!m��6h%�^H��`��Q�'"��Z�� ���'u]��Tn+6p��S���ev�c�W�RJ}�J0�@�_�