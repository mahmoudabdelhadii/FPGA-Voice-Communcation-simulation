��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��,�y�}�ǰ�=4d�H���`I"��W�`r���T:tB�T4D�m�)�	1��I�t��
��8(�8t>s)ו�."[�漆���]�~�]��;�O(1#5�-� 偙O��QZ��~rL'�x[�i,mׇp���O�I43��4d�,�H�����SN��d���3���r��m���̨T�I;uj2Y� Er�*p�Q$Gm���p�V�`�2^���,hz�<p��l�Bxt�5��s��\yq���#�@W���f:m��T�	,*�񞭋����_��㧋l�	�\�:��uGd��PǷ��N�I��_����Tuv� ���us�(H�~�{2H�:Zor�Q	#%�3ˠ!��iS��95�,?�.���/�F�i{#���Tp5����Ҥ0{%���2vpn���X�����@l����3dc�ק�3	�Ed&3�ZN O���z��s�yxӡt��v*}ԫy nj#��lc��m戭k[��5)�A#�����8�!�]�Z�s�M���t��w�!��'ÒE�rv��Ϝ�c@<U��\tq+��&|�&X1)C�����r�A~��B�&�����s�:n{p��͠R�X⺂L^��R����c���f��J^?��ܣR�O 1�rV���:��T�4���AD����˩�F�w��)Dm�O�b,�a���1$��c��7t[i2>�ޔ0,S���󧇳Ϟ�ᒨ�-��}�!6��Jyv�醊�^_�(�H�(y^����o#����X��3-�k\8�M�T�"`R�DF6ȕ� �,5�;Ҭ C�k���1\������k�t־9�}���� ���QHF��"��t�9 ?��{E_�7��!����]Zɬf(�'4�o^d5��o5�V+�����YE�٘tv~ұNVz��!#:�C������w4���}�A�X�a�h��2�),��ۨ�[�s9\�^��p�%7�
�L�ƕ�9^�n%=�)�)�NB���	[��w�o��9����f�x�\���E���F'�Ɩ���g�5�+�$
�H��6�p�?�b�O����e���������z�w�?�������j)T���T�\L��8y��=�~���U�Ea����r�2�Ҿ�+4��^ȻI�v��d����{樂�-�l"��mj��R�)j[��t��D��ds�����mh�M�����%���f�)����.�Q�aBR���r�v������JYD˨6�LA+��x|���k�j
q|�g��].��焟�܆?�3kM�������눋�r����?5i��j��Hy�N�|���}�tɚ��0�|SE8/O��t���JEY|�Pd�߯}�����4Q������`�_�1�oe�-�E����L�{F�iȘ��X�G����r���U��)����3�҆�:ɵ�
̴X_e�� ho�"�΀'�c� ��=l�� Sw47��7�a��}���,?�/?A�84J���>��ֆ�>O��=��n�`�(�j�7�-f@��|��q��}@��AͯR��^��� �����m���s���Uj�֍��rX�o��3��8I��S!�E6Ǝ%�����P&H|z(�X�J���H�.X ��&c����=��?�����=��#~���|x��C']@���cE�9����ܝB�(�9BEth1�T{Q$�<x��,��v����D"�QDݶ�GT��&Iӹ��F^Uܢ�!�U7vշ�J���oH�=�b;W^�Y����� �n$��5@v^7���3�#���ym{��<o�r�˷�P��,"���M-o�w���$��_?$6䮭�.�� ;g��E�t��\y���Mr8�mh �ӆ+B�u�yת�c)�ڦX���x���`���A�p���J����P�H�נſ��$ט�:�Q9���&���>G������Be.e�`uЉ�-7bD�N����b��!���cz��o��؁B���S�y�9x�+{p�I��>`�d��_,��+K>L}�(��QHX��ؔ]'�xKT'P�'K�<+���oO۠���
�pi&����턴��R{���T���l�{n�ƀ������W�gٴ��1�Vj@X��{N���,c{Ũ��4��=_ݽ喸%\��wu3-��\ X���P�ܖߪ���`�<�񴭲���4P��T��$l��l� �ϔ�af6橖C��ab%c�U%ғ]��p�Gj��i_����?cX>�#���+_���()��(��tO�KM:hV>Q��F���|�b��bE���6A]zg��(L�d�.������n�8<�y
��ӷ���8 +�Df���������q���R�����h��;6Q��@-;L2(�v���Tq
�L���7q��<��Y<��2�}����Q-�/��n!�զ�H8��� 7�D�Ϣ���<ϫ�� ���)�z�~�.�!$�j^.�q^ͭ77�����p/ZI+�J_�iyY�Y��$�J����a�W�RZ�pq�\g��U�t� �U�e>@��F"T�{��W�7�st# �m��Y�+��{κ\�Da���oi�@���}φ�<��o	��&��f�u�羅���c{?1`�E�&�<�7�I�h��t����%.ܴ�2���Zb�\Ya�<��t2p������|���;�{�����?l�[������Lq�bֵ��u�M&?��-��'�c����}4������H���~3��x����v8+�	��~+�H�U�o��HP�46=Z�{�������,:{z��5�[}.��*!$E�>�tc�W��=� ���G:)Q/�Bňڦ~�B̔��dΩKQ�MF�>����X�U�8�n��%�+v���~�h/;�av<�qC���lK��=6"���{zRPx�+�-��8�f�+��y�qA�/��*��w����R\�^-ؕ@x��rMV��(������
R��$=��9�Q���z��=��Ցc�^J�A8�?��de\�Ƨ/g�E��#�M��8��V!�=��M|-.(�-��V������c0�Q#��瀯S)Jj�1K}�pG�U7��vø!m�����q]
��� ��ZgƟ�z,���e�"p�/�34�����4�R��&`򿸖B�:�^��ާ8
�׿�v|:���fl���eq����E�(�-I5�� �LX��xs���$z2Y&�Cg�t��B���ݐm ��ȯ'6��W��>����l8��Y��NE���"�k��ak����$���ԁ�p7vW�;���q�����&q=��}�E����bQ{��N��;V���#e�qQ�*g���T�ek�M��i��~������*5�m"B��B#`�)�8���a�`�󝂠�XJ�����_��-����U�8���!<�3T�##�;�w�zd\�H�`!���DV��n)�-��%��g܆�}׋�PZ|�Aj��(�'B]�,~���}D�WV�[���@>���R��x�?N�j"��S�c�#�6{}b�����B���Z�T�xGFi"���	�P.�i���� �܆�O|����E�yaT���
u �ս���s���B��ۼ�r�����E+��A�5��0�*`��Z�D�Z?Y]^���p��f���z�l����a"��� �<Z~�
a���ރO%wJ��/�p�_��ڕ�6��=�� �1���5$Bn����� ����$�U�����-�!�OTӃ{.��6�-��6�D�ihj��T����ᘽ$<{\�9�������GD�YAG2�.��tJ��Hy����=ye�nS0��1�V",��ܦ�cʥ%
��>��415����iK�-Y�$�f+�:	��p:\�)�{O��,��ޣ�;��u��#��,/&yh9��K(�w�}����:��t��+�;�*tբ1����gWfd�b����'�Og�n�hT]�t�j�_�TRyb`��d{v���ƨzsJ�hX�_EpD�M1}|��3di��^FR���L��Yxuv5g��T灓���FW�����i.�Q^��}>dr^M&_`?�
�S����ƥ`���u��Q*(�B���ۯ�\�s�4B�朢�����"��P���!v;1�Dbl�!��V��4�_G�cv<��M~	A�%�Br�.@�� �T`�3���$�֜z�_������!���	[�����Ѐ@����F6��J��׏6GLD����4�&S��^gY�����r���Hhw�Ɗ�5�$��S��[\��d���6�����!h����c0DPM�g�9�Zq��=���I4/�X.͓\x�0���`�ڼR��z.�̩2��,��%�8m�?dU������#��H"T�FD%ǣ@c{��*�����B�"c�E��M$~�TG
opo������@YL��&�-e��)�['O�on�ǘElx��zr�j�[��$�847�b�.�`ȆHP�R����.�pқ{=�fȲ�mo�_U��<���z�kV����H����6�E�RݏO96g�u�K��df�N�Je�b�F����F��~A�p������.@[�7S���K�z(��앬���	��	�!a6�-�,I%e��zcoN�v���ח�gl�؏`�M¥�P��5�O��/��~Z�
	J�:w��]�\�ߑ����X�8�w����<�������j2�$��~���
p���'�+�6ۑz���=9H.;�8�Ȓ)٪E�]��%�}�.�AP 0� 8͖���n�:���l�6�㯓�!��x� (��ık�1'���%{��E��ё�;�_��fOf	�E��Eh�g�9t�%#�{�Ϧ�O}�Hw���:Mi�c�jR��?�K[�5�O/��H�x����"���u��;��d�Ɯ�Tm�]10,��-dv$��U�%>�a)e�X��\k�/>KK��QcY�#מ��F��4��5H@A8՗�/�vu`��fb��`Y�K/��������x=-�9���z�4񬹳Y������(�03��t�UѢK;�-{�SAv���H��u�B#.QkJZ�b��b\7�RU��g��̟	�[�	vr��M;\�ӳl�v��$����^bֵ�R&[/��8�#��(}��wx�܃4Ҋ7j��/tSǧJ�Q�yl�^����v�>�`�o@;�-��}�CF��V6�����n��'C�e퍉�����ȵm�᳆�F���U�x�b��\kt�=)��:��p�0�R���C���z��%����3��8�n��!�m��p6�d�6q�����k���Kquӽ��:��]��]?E���ҝ~$���U���ͥL�|�n��Г:b�j��x}� ��:�#�օ��#}�N��*2��0�N��	G�0y1�U%Ns��1h��pȺ�� �H,�����2�G]�:����%�_F�-�a@S��Mt$�ٿ�{/����������0鮆�flַR�	�Y��������f|e��A+y��t~�߸�Ny�q\B��+)+��Ĳr�{�T��5�m����\4A϶�Vm�{��l�H�$��A�y�V��Q2�4/s���X����,e7��t����z�:�u�C��#�+(�M�>F