-- (C) 2001-2016 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
KEv+PQZmJWY4JiMadd0pRtq5mcR3p/9+NWTGybb2c6OU7sAH0vaAEJzihkoKkezeFGDyyHIHr3WI
RUWyHyblAnjkMiRG/MG5e6dVpG2zgMYr4DL536NWRbVkzFxVIRApBzXRo178HZBzFZf8pGABYJrP
i5CYBJlqEkXfBrs6k0092JfgiZVD2fgTAcLCaGB5Nse4QUarOERpq028SdRFXCz5IrezaFbSO39/
e1ouXF0WX4iqCGUW0rC4DYHzIqmzoTbTeV3lTXtowP09ifujH4k/meU8RCJb40fRpS1BXMDRIUGr
U/+HSkJtv25PKeikhBCs2ERkQRu5VPiIXwCvHw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 5184)
`protect data_block
fgjngxRGEDvBrrOzDlMv1AnltYHqud7CArumaSrGVMrMzig9fDyCicnla1w0tAanASblWLWYZPaW
w2rLf+RfOMnC99mwdJIGN7kmi5cxmMSGXHkMnHC9mDe0OfDCSA0CWmnqrDIEPWQJFgcSqHkpJV8S
SfSPFKhgehA6m5agLzOA4yTPFyqjR7lP5P0RUWGesXEoi+IC8iDk32e89yYrr8pedRP9WEv8ANx/
9Ue16fZKnj3b7UXM/tscxrAp54GBQtfN2UEespAFMbZiMHGlEWQy2kBspNGBjajv6PGBFindFOhA
xybQPDfQRWrKkPz0IJp7N7y2IjyRSbWiigIEu/0orSbqek9A/TU7uKc8EMSq68AAAPOkh6q/Niit
GpJwH48Y9Gaa9Rugq2Iwhh427vh2s8YcU7QeBWsJ610r4BT5D0pAZ37fb8YBl5Cp2gdvji2N8VuJ
r8NYkOacn0bxyPhweB92sKDSnbCJ9+r1BCzlVposu+33CgcB6Dqu65fmjsJ/dg4xeye+htgMp/Pi
zktWME9EXgj4+LNn8NBRiakjIotc2JpZU6hR1BbuYQdCOwrG/Ar9ncsqNmT9EeVx6+ons/8CifEq
OmImMhYegMQuaW/Wh25n8/Ji1Wjf30MNBCCn9/cGiOtuZRxAw+efMSldNTYwTz3XW/jQOQsYs3d4
uOqYAPbSx/2ozaflqBTOs1+35XWWTqvgUlsDeCOtGQ/Qvuk9cql8FhxacRTEhm1DiE40vGqHDQxu
9FwR+uL2x68jyujX0pddjh2Ta3Were0pNWgHNARG/91RTDKGz7R20wy9ccdxhFc2auJWeyGljlkD
YTTczQXIifTE0p4hGjuiVYg3pb4GU6MwntsY1dhdm1ApDbsGslbwhJN557/wKgFVmCh5WusvrXJl
IFVfDcJ6zw720eO1w6babh1kp958GIBPv1ki+DC1XZWyW2ECDvxLsjF0wphuqwqkwewrWoVHNnCR
xx0OdopocAg7HtnYnwIEe+Vv4Kjsn4wW0FCTRdf9QIV3t7VxCXH2QOlu31HxDJTQo6r2OQhaMfJn
3R8nqIktWxpF5F7yc3uRpheGlH+w6XkOP0fcD+93Jz2fo2I1Ee9wCH3cchh8bgF0Zyeuk59lNa8Y
FvwNPgvkNbQNYgUdrs2Ki8eBzoDCAJG0YB+e/HLWH1cKsMRNuqhvTt86ZEcBSfa0zrNV8WQXHMwd
zN4rmiJPfvDy8OyjHckBfPAFROMOpTlyr7+gc5Np3/TwfZ5P+ezKN3h2rDmeIFymqnu7L0xXwjR+
wthFJMUgA0Rsw9dweL19UYNe8Vm7nqfF2Jt9hp/arbD/VSs8GT+HtbcFN0NT0kiRXOEAkoZMsOXd
VhfAZPrNpuhoadv67ZRB1vhxqsNjA6yylbh6mESz1c388vD8BXzuPoraqfOr3mVFQpbl1//4Q/d5
ryIBOvdq1j2dlUt6zQmQnVgg1oTbKo4+3fQG0UmeW98q+p29+50ZqoePu0YgkLusMCOq1MvR7iDg
WkuuGBfqWC5x0lpq33mTH82Sb8HAhDikaw31KxlmH3a6p0Ma70zuigj44jcMdMJfVfQ38FxMrTK5
14ZxOKoAhrYgIvA52mxvx5Mb2xpQNCS3kr5QoCrLLyRz7J9TMmnLAo0X66iOeYzQA9G8X1d5PZss
nBp5WdCt2t5xWnbYYP/Cp9xFx/jN3uGayQw2tUQoIuiMr4ZdJ1aVfeEd42/qLWByxx3IXlAOyoHR
rGv1FtVvCg+E6cCIs3kQOi0SU8GLyAKniRGnFioN11MRLWlbV2SvMc4dmrdH02khLaRazpa8UNob
EG6YxSVn0LjyONXvgNEkgaSGEa/g/e2Ok1/uLnp65pXYIQQO9eOOOHjT5FAciis40GgxkD2ryEBT
CAIAAljgrDSrs4xK5el6EP4q4tL23pUMxrRn1j9eV2KEj6vc06RUpTPPyVmWRWlsHRePO5ZoINzS
kn/VHo8qR8eHQVTFiyWQNeegqdBKgaLyw/3IYutabIBsZpgz/praEYGL+AJMCy4GXOZjCwLHzmjL
VLlmnFi07mRqiO+y7eSQFLCYzUP21X9s4geU5jNr8Sj5Tri+T7bhOPCW1pQKLCXJcx8LQ2puIYfN
uXipoF8AFMFa6A4x2Z8YEGuFpm2npAJG7uQdTJbyGEBCNqiEmkzqXDsW2rwDZJRc2NWQ57WzElES
ZNo6lvgRK/KUcQQuX3F3YW+gkkrYMol31oTTIM3k5umJi1ySRPkAtdrrRvAJ0GTF8Vt/ldifM5l2
8EKkBVHlRJX01fhcWv6lGhES+UlA0kWtSlhapFbFU6vvH63sOq32JyTg6qsV5waga6Xfk2pG6JSM
Gjs3h/kcmkPIHNOHsXqPWFqwqHgklh+C6bdrggygFnSfrYduFRh8z/+H86K79+butu6ICNYhVIs4
rmmjt3fLVA5yvVONFjB3Oa8b14zANDsKDUBLBf5Hhu1AIWaj4YHMsxQp9BKw425ld0wzvIjwhVan
TnmrVUZq+F0+hZlnbOjBkP0ErFyi14ZO3E0GW8+SEq0nUULhIGgksr8MgyPYnV5L2B6jQVhYgJPe
mUsfXRCltAGmj4czVzbdwhtZvqixmjOhwWgTiTnVuEVK0woL1yqREPscXGnf7RIh0gtEZKw6/hmY
1wRcQKDHf+sXyv0AI0boqSHln3d7yVguAyEcaAkjBbaU8yXZsPLpfmJuQOV719W89EmHLYSaauYb
o11ZTLY/aHuMhlp8vl0Q9NGXrMcxga3sncPBEewCpSbMu6L8s65IG1VVp0uL/iT0+MFGtye30XTe
ijEHMs6IGe0ORjPS1/SWhS9BdaiAFiKG5MEXvNDHxAmW2hJy1ewUW15eJwbX+CRThFcyfEyJif6d
SwPor89nBEBUnPJfbX6zqqx076l/DVG3J90k1p+gK4wO2BQpehn+QSImN4thLU3oQjIfsHhpHTH4
zR/b+nPL5FlVqQylnR35zT0qQKDiLxOJaSrjxFSX2TQmm4EkjqpG+C07ZLsDmtzBPWjAhPYs0mcH
xjo/0Fbcu4R5vkZb5P9vju4a6E8EjLh9apq0oDGFqhHdGRCGKrtrTxmK7CRO/WEdD9UIGIqmqE+B
vcADg5W3LWqvNqaFOZYn82hblElxyTr8Fm/ToN9sQwtTqSQe2UcUft9jykOXN2+gjkSBlrQk8/N4
tmuaBGnLITRwezoZ81GYj4/tAYh9YozSBa6tZY956r/V2Yo7g2jvgp4X904W4MIZLRR0pDu6/jUY
J+LZy7t0GkXq166GQlB2sQhBBPlgrU0gIMsmQJWzWtw4YcS4BZ/qfRPNtVkgyt9ujHy8CDp1x+bT
1pLcWReUzwGUohblKdIb4+8XrBD1NjHx70pOOZFOEGH5G+XCn5wYdztR9+50f5jIj08kmHy0vuRz
orDR9d8tthWckkxWhZ3NoF7KwLCcERadl8SBSnGdb1jMiBhR1zboVxBNy+V5xN7t7gsWQ+gZxZ5H
7iVi6kZssNldb84cxKoL0k8xCHGsc0OdJCs02PhBBpa3sCQqDJyZ/EazcehKU+Euw7lHU1IJqpM8
DiFNYclxnNQ35n2wbh9alpmYGM2fEKFhuIF2/0PLeIB1wGINWgCn05c2aIgGpbkhExwZGhG2yaqV
gEBspIpTdxGLlLq2dzjDZeUExCpnNx/1hfCWcs7S2xNiBQ/GJD9zE3MIn1OB8K8VUtbIaecUkh7o
Gobs1+a/I5uS4J87JCOvzNAiBeFo00NJuCQBewK7JQnGetODxh0rnThcXd0E3pgwr1kgyM2qGDdq
l5tI9mdS00tV6zkRNoTU0kB52YCwhQB0V2se1ukvYK/G+IyRAR+X+OmCuks8g7aIXI0KyxLm+2Fk
xIW5nMfsuZl4Latknnlwgr/foqPmnGf8fkcJr4aiB2pFOzYMKjF6hYpzU3m1Lz0BNKPdLE4iAkkp
JvOmMOCfdW3yUDauP4uiDvbbGXGE1LYyDinVK9kYw4W2oTRu9qYdyN//DhwaxQbJyGxoZc9/i8l2
yNlxurQf61j8dbe4YADcj0Vdn25Rsp11IFkpf0kp/R4TchnFEbD5sf4s1UoXb3yRR0fOrvNTDJwt
q/wvPAvZIMR49k9brRv4XuQMGbF9NcrJK8ORsAKsS/2Vo5J42NsXO3MQgXQXYILGlKUE8SyMqq2b
JEiUCT7uhyT3ttJ2IpeSC0tYAArsl++qMljC769P3dxqJJDqHs13pzuLkvokz9NCbwbfeONCejjA
OXvnMtScQ8PXBEJMOgEj6acuB01BLutX7Ww+zEZNz+ZoA+HKU5aBakq5lihtjeMOfXPuZ9xUzdDX
ZZNgYSJA2KDWKQ/5tI41BVrxjgW3ljf4fVhAw/8/UnGPvaUj1maBkmWkoFKY3LdEp09HZ9QVsyqx
5pl0kTY6V0Aawm2WP40HvxUOLyTEBiBL28BEinJ06BdH6sKSJZsOMmL9zHQBwOu73SbNB4VSpsX5
CN/Mr1LRk/QcHqtBcyXdV/uDbstT5sh2p0i2O4ivpELSJ5AapAjA+Erp93qcPVN0L2qQeuXfZctG
Z4MdUvT6JrcSc31f9hcdywBxcQjZS7EhcIAlaQ1oh5TpH4CNgfuWKgoeDjSe1QxSvx5pnBDyTGmN
WMVVKvkjFww19tYte68ZTLUI5yzFpJNShb2bN8ku5ttnmTzZSF844YuggYaUUAb+xpTqBYSxCTb5
fs963Gp5CV0iw5LoUNibIEQ9mArZDfqD1R60gx/KK1G9cycfnrq401s3WP2aZuxV4SUyi539RZcM
fnTHLvYqC770ccZnE8ekGAk7QEtZ2aEQqwBRHVzIcNRM64NVeGKv5sbnB22b8K11xaadblRiU9qM
MkwxsRvmjYEOqVst7s1uicMjO/yJjqbxMQJDCctmRwWG54RqRVyTwmEjRffbvvqXUYE7x4WA6hiH
MtEXUBp8vH60gf+uOGzQqBJ9huL5wwhmXqYnVSPGckpUQSsIpNchsogn6UpymIT54zV/Cgc7S1AF
YZplL60Zl0EoWupeikzmh9qyVcbuvG2jSuWjOqxOUw5XHFKx7iNx3thHXCBStQK5kw5P8HswlP80
qFG+lcAQOo+YMN2rzZViuqK4dqAHo+UMUs329597lAnQ7hb6FIMqCB6LhvfFL4YdW7uy6knjmows
qyrHa8TuNeb6yDQQ9E72jT+9ahIGIB/fhM5v2e+i1mJJroKyI93ye+BvAay4y3BqwjHmpd8j17BG
M22jay6YmALc+OmqCU6atOQHHFwPTREZbeqVe8SyjRQrim78ZRRThRIEUG9kTvDPM5rFBC6B0m8p
NUQzRwMPcB8A26ijwaoNiw+7+4gQZA4mg9ChNb5xXwKc9+Dor/1I6f9e3LmgGHftDtqBOMC4u6mt
aJRcrYAirpQgLoDpqYMVNt+COOZFmw55PpKsVwuIislMFcahhlikS61U2MT7njG81ouTE2ciR11J
Xg6zI01+9fXw6uOT00WgfyVS99ejXMod9NkBmJJT9/KowJVPiMSZXLs5i9f9ZIT8Pnq5+V4KVjVp
n3+pEBGxRRiYjn7CNOC++fpmlQtRN0eFd3wmz5z1+Ta/7+dyZI2gaAkjUEPHqf0ziaC0k8o4c46m
iqKdXCeOd3z9gFf6klvLB6d+ykmT4qqG8ijU4Yke9ek4nHD2X19CyVTJsoP1+gOki2VBAUSdUDN8
LKA32zlUQWkkAn08DfKhiVaTla18qGmLuZYSf8hBnrT9ibe/z91nt3jJ8kl6Kcew7453sO5w+Sfh
1Ft+dXPSTohroDcH3Krb3h7JLwxx6hrytdsloWOf+c7tHDUjLPx+MkOIpsbBB7SPOgzHlH1if/fR
dS9ZcpW0Cb1iQMgK7PDzbckhqV5gur0mdppHNr1/slHlSULczOsGmn1As+ccj5W6RUJ4ixrY/PEO
VOiC+MORQlepApALRMapsvqr86WwF9ylAtHy88Kynghw1WiuzfkRdhbZ1VVwFxTClqvmgaUBwdYh
jXI0hxcZJxpRMX71gUdF76NDSgeXFY/9DiI3sm4nmdP7JbQWNw0HuchzUpQjCRMYokOjTOYWOSsV
o2fL8HZV0nggrpoWJddr3GdG15tpxP3V8AqXkyy9+G9ncB2gpeKQKt0KjCyxbrpOfgB21VB+QvIb
NW54yeUx6VxWgmq0/VfPSe1scC4m5p9Gx+ukeHg6S8k4Um/uTauSjPM0odsxiM2tIv+zXScuK1CD
EGt/+hAfCkp3OL1f3Lz0VsnU2st3HBBaXCaKkECskFlGvY3vrDgS58GKQ2vRweAtLNVFhh7wncVR
t3C6Dd1fQno3tu0o+FtDWeoTJ1Ku549Sa7fpCoSWy858hXsx4H+DMyuSB4SAch2kTC3fn2Udx7K0
7r97hfLHSdkCeBA1hqSRb+daqeivqWeXNsjrnYrHtt0+HSz9zPNTXTQZeNcSGh31OgMoe+lAdZTv
XB7MzP8tVI56xLiEvjM3MGIJaAChEwGRkuXO6xYPoKGiyQDFPnP9u9S6qdVDFEINR7ybrKilwtF5
FaC5izBm3cLTUCnRSIiOHUzF+/gAqdXkCty9OdG6wwCL2RTkJLxSS/pPuujT3ENbyZCyDo8pYYQj
mZTDlW2fJsJEVx4vRiOEweqtr/93m+AtvU0vKgcZZPlaOzoZhoED8UHkAUaTBR4QOOCk5LsmtZuP
2uj6Vhd3iwMXXnhsLSnXC899+1WTUpO0Mp3viEEgvTJThpP9ox0EMnUYt5k5gjbBLkP5KpHme25y
kxqNk1FxL5CI7DsDSbLmgRU+JjOg+2zm9jm8P+k8z/zWx9cteK6ELpzJ09hi7EDKPrFf7/D4+23B
wPsj7soBZ27V4uJGILvq+07fE8ai8gZf8Nodgv6t9WqfMopfIwB4XZGU7LGolyvG1/RqhAXb
`protect end_protected
