��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����N~@#�k�0!����+��=L���0�ԴZ�2�Mc���ZO�����=�����վ�	"cqw��a��TS[��{=:�����K��-�մ�(��k��N�-� 偙O��QZ��~rL'�x[�i,mׇp���O�I43��4d�,�H�����SN��d���3���r��m���̨T�I;uj2Y� Er�*p�Q$Gm���p�V�`�2^���,hz�<p��l�Bxt�5��s��\yq���#�@W���f:m��T�	,*�񞭋����_��㧋l�	�\�:��uGd��PǷ��N�I��_����Tuv� ���us�(H�~�{2H�:Zor�Q	#%�3ˠ!��iS��95�,?�.���/�F�i{#���Tp5����Ҥ0{%���2vpn���X�����@l����3dc�ק�3	�Ed&3�ZN O���z��s�yxӡt��v*}ԫy nj#��lc��m戭k[��5)�A#�����8�!�]�Z�s�M���t��w�!��'ÒE�rv��Ϝ�c@<U��\tq+��&|�&X1)C�����r�A~��B�&�����s�:n{p��͠R�X⺂L^��R����c���f��J^?��ܣR�O 1�rV���:��T�4���AD����˩�F�w��)Dm�O�b,�a���1$��c��7t[i2>�ޔ0,S���󧇳Ϟ�ᒨ�-��}�!6��Jyv�醊�^_�(�H�(y^����o#����X��3-�k\8�M�T�"`R�DF6ȕ� �,5�;Ҭ C�k���1\������k�t־9�}���� ���QHF��"��t�9 ?��{E_�7��!����](�S��0�q��w�9��=�i]�1�GʦȪc�W�XC�|�$��}q�6�\�\���Bp��~�1��<ΐ�%{�%�3e��)6��I�*�K�X��q����y�>��sR��u2��V>曛�aŃ����Ur`iB��O���b���	�g���<�%>�N	��6��1��h,�f�׿ϮU���C��@�\��`w��`�7�L�'Κ,�G���}{3�1�g�?�,����;6�[?�+�pI��-�6���DXT�m� 

�.��I����	t��6�Q{����j����mr�̘��9)�5�!qgo���'n�pK���G��B�G5TJH����U.L�Ǩ�	Ɓm��i
!:��սl��7�].����Tė�0y�P�0lD@x���w�|���A���dA�y�l6SIF��gi�8@���$�L��+w�/����T�%��S��fq�|��
�0��%j�(��l��g&e��4cOճf��%w�����n�f�AH?����*d��� �Ϫ���q�.�4ُ1K$����ܾ�c��t����->�A���6?�✱`���U<�H�J�qPG���B�S��4<O�l�����B;{=@}]<'I)9�ض!����O�[�St��a�C�˝p�̙M�T�|��K2{������U"k��Q�-sL�Ӧ���	�����e|����)KY�d{��v��䄜@`�X%�����!U+H�0m�O�6��$
�"yc���uM���VV�������&�>~����s�S �S�-����L�0��|���ڤ��w��ήvܣ%��G��W�n)��85
l�08���)V�*d��B���y�������=���y�%���65C �l]�D ����.�9v&N\&��P��/�ϴZ���heI����solN&��j�E�	0F�g���#⬭`@��}h?w��Ȫ�n����b��FrK0eJa��+��:���C>�u��zi��K�u�1X�܍[�0�6V�l�y�������PM��Ɩ◅��l��H���*g���ju�F��W�&�bi=�D���#s)0�~_}n�¢_���u����y�J�|ynA7��Ʊ	��Ha#Kαz�1�h
!7�GM"q@�S2��_cii�m���G��悰隸Ը�<4K�(rA"��W��)��ʃ>�G,��?��Rj�w;n��qc�ㇼ��+s��xs� 	�?`1���#���ҽ���Y�mKk
�{-xVE�X�bS!��ugMh��D6��� ��#�K�	�t3�a|IuB���U$���'�����&Tӻ��~�oOXoIܡd�`^������J��0|+�n�_|�����Xc�!G�*U��2�J�!�?	�B�2�\��z���]���`z��p��.�ķ���S��P��6i���L:��@xW�hʣ����b��̋Y>����CbT���w��!ΛZ�Z�!�:�{��f�x�(�e�	H`����Z~�H�����_��$���A��Y�����L3���D&��K�X e\���5QI���qb�;?T���sE��O�c����o��t����e�
S��p�x��k'C�y�z@P��/%d룧���R��!3_��?fʦ�<���מ"���-]��<���5�pQ��;E��E�Q��Y|��u0���nWr�s�d�w�U Ek*����g���Wkӹ�;2$��Ec�x�C�y˼��;<?I�c�L �&[�;�R_���{��΀kQ��0�;S���y(	���|I�sl�\��Bh;�Ck��h �Mc�o&̾�!oTo�j;c�%פ�.��Q��S�G݌r�yz���k�^�ގ���q(�C�B���7eQ�^����ʹ�,�-����V��;�u�$��*����9�!���L���&��[�dvyd�L� ���Ɛmj�*̌H���{S�VŨ�9�⪿��1����m��,�aj�Y{�v6f�T��oʹ�OD�@�k�1�4��"�kN X���w����'g O��AȽ���^�5-�����qM�l!e��׾�F͒]7#��i�XX:�@��	�yS��P�\��N��_��Vj���H��C�O��NW���s�(zWHA��P\��<5o0����"��-p ����n�ˮ��A�O󋸇�l���ǳ�
L�M=�X^R9��?9��H��:wY��6if�H� ���e\��a^�wuذo�_��'��z�m�w�4'8}�ġT�U�$ٻ��`I��ume2��b[D͖N�\@��8!'��9[eG�Ψ�_{�3�E�qFl.�@�lK��|�ʍ%n�@f���(�'��wkjh9D'�`�0!����D�M�@�j�Qd��|2B�2}0��70�Kvgdoq����t�C�0K��{�#�&��ʳ(Sl���?��Z�Eպ	��ۼ�Zv�����'bd�v![������P>A2JY���.���j���7߱�%��͔�䂢��ٟNi��֘]�v�G��/%��3s�r��g8��a��o�k�sx�B�Q
z�֠�:�F��ǐvi�ij�P0��$����
�}{�w�#,w�t��������-�"��"2��N1���LQS���R��R��I��P�g���ZT��9�T\\��`����hu�N(�~gP���e�0 �6+
I���v�ĩϻ��
p�^=7�E:#Ci�\����Y��X�T�a�v3w��]�"�>�|t6�.1���EJ@�"�B����1/|l�/fVO�H�d��jsV��j�}�zkYf�4��A����6��ݑ�%�aFZ`$K��Di=�)�_�/�"}&	-*&�V��;jy�ݮl����;X����+�ʬ}7�G�����%��#&�
���x�fɺg��49~���<��3U+A/d�џ~R���V���u����Ȋ�8��&��:�G@c�I+ ��u0SI�*�*������-�3γ���\v�j�3i���U�_�-S�[�"s�	�Z�gN�q���T]��x}y�� �k�^�*�V8�R��璴 v��/ap�u^���@�6_��mgR�ۋ��������[��Q�-Q��s�+�[�LM�ߛ�j��aD�K���$��<��i�X|�l~�����´���ң8m���8�P�@&��%��Q��p��;�������?#�K�(�u[�T%g9*\�4���W�]��\�Vj��J�c?=�Tm����
�M������̏z���0���+_ �R"�,Q�P����:� !�~�?ŤՇ,��l����e)���w��N�t���^�M�'�el��?PNPA�M;��������8���
�C8dݱ��lf���%��σ#`�^:�漚��S��+���fR�����K�x��+hhy��&\��M۔�;��i���/���]W��>���}(�����}��n,K��4��wF�|�v(��S50�E�ᧁ�￠�P�{ph	jc#2�I�����x�s�?٨�aO�w���&=��>������ˠ��:�$\Y#�����u�X�����I�2���=��1NZ�[]r�ir�*��,�na	4�P�u䁪�w���&~/��?��B�߁�.�5�|����1��R�s��%*m�x��H��n��o�P�
�b2�5t���]d��CWc�!��ÿ#G���ya96�v�A@!����jy$�aj�o��^�빙O4�q@��O�EX�r�J�/��9���5w���x���C�g��7���/	`abs�����K���K�ǹlM=R�U_��r@���	��.���p0�_������z>ĺK�-��n��ܫ��1y�m�e�_ھA�/�^3�&�!c��V8W�S��Y��5�f�������!���z��=Fw�Z��.�;Ya�OWƨ�!�[��ʚ�ѴE�����U��;?W��Vk_�-[e5�F�n��Y�I��X����1Z�+9� �E��ɶ�#�bݴO/�B.B�Wʢ���aE��D}upW��
����Uj�ڄ�����ᡋ@YDD�|�}>i��q%���3�FY8Y�I�K�2F��i4\���:�|>�HI7�-:+M��{�y�AE5L�f�<��;��Cbp��71m�ｶͻ�ǔq
��B8�s!��G���Y��}�c6-��Ru�������0MvhS7��#�)��%�h�cb:Ja��,)^Ź/%��͡dZ@=�^Hd��N7�/�rmY��nA�����C�X%8WtAF�0�ptF�F9
��ل�̭i3���ِZ�8豳;le����o��9�����
��J�-_��~�g�Ńe��J�����,s��Wvk���u�����U[�0�7���L��x_��U��qփ��+]Z^0��ad$�h��Jp8��X�D~ȬJ��Y�`��G�X����{S{��b�gD�ao�����Q;���l{��^K������o�����S	���O�ɱ\�Y��:mƱ��l^LjH�_ �q��&$�.�KD��01��"�VWa_W�s�G�p[V���y'/6SQ��T�0ω���ӂ֤bC�VĖ�?@���aږ`O�40B0��Ik�l9`P��k>���wr5R��mD���p���0��X�ٕ~B	L+:�)Q�;Ĕ2��W�)倕.��$/�3������]�3�啾�p/#�Ҝ�@.ߧpf�kr��e�`}�)�����a{�F����,�	���]�3��Ώ�i�2���L���$��jҐ�Q�W'M�E�(�>[���L���ֺ���������-�ma��G�O����Y��	�&2M�p\>gU���l���xwW$"�_�Z�}c3�C�G'��Xd.ޔ��rm�Jt7ӓU�����8X՚�#�-���3 ��ǰ�ªF�7J����;�4h���g'�i��I��u#��,r!�c�s��Ç��8��f;�եp��9 �W5�:9r���.f���ܨZfs�ܿ��إ���[�$N�߮�`�gx�c/�A�efǭ,������;>n�g׃�Yg�qK��b�������#갨�h�v���;��I��#?X3g(��	^Ȩ�Q��p�|�j���od�8
kJ�sv{��a�lz�,F8�ͰC}�?)\�s<�!ܫ�hϙ\ƙPaV�������$p��mr��#�CY��yS�����M. ���&$p^+H�Sm�Z����L�wY>�~�Z�_�Ѿz?Z���(����NYd�їk` �9r�確�
�*�=�=���XvU�=���|�KWE��O�~��_�O������Bs)�Y�~v�w��z�C��Vc{��������iә��C��g��_�N.S�����>w��K��>�J�!
��)5 �W\v��i� A�dj�
�X�7c;�j����L�؏"�6ʄb�^ê䉦��|Na(�����G'�n* 8%����Z	(O^Yܵ�"ҍB�em�F����=*�9���nT=X�V�$)�j��!r|Z �LUCYP)���+� )M���&"�w�ጿ���Y\X:'9��c2u_��װ������Wԙ>��eD���	���X��:�(唘�HɼTO�O[�:�������u�5HU&�Nb㈵����C�S{ws*=>����