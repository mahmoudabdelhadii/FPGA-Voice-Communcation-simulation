��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��,�y�}�ǰ�=4d�H���`I"��W�`r���T:tB�T4D�m�)�	1��I�t��
��8(�8t>s)ו�."[�漆���]�~�]��;�O(1#5�-� 偙O��QZ��~rL'�x[�i,mׇp���O�I43��4d�,�H�����SN��d���3���r��m���̨T�I;uj2Y� Er�*p�Q$Gm���p�V�`�2^���,hz�<p��l�Bxt�5��s��\yq���#�@W���f:m��T�	,*�񞭋����_��㧋l�	�\�:��uGd��PǷ��N�I��_����Tuv� ���us�(H�~�{2H�:Zor�Q	#%�3ˠ!��iS��95�,?�.���/�F�i{#���Tp5����Ҥ0{%���2vpn���X�����@l����3dc�ק�3	�Ed&3�ZN O���z��s�yxӡt��v*}ԫy nj#��lc��m戭k[��5)�A#�����8�!�]�Z�s�M���t��w�!��'ÒE�rv��Ϝ�c@<U��\tq+��&|�&X1)C�����r�A~��B�&�����s�:n{p��͠R�X⺂L^��R����c���f��J^?��ܣR�O 1�rV���:��T�4���AD����˩�F�w��)Dm�O�b,�a���1$��c��7t[i2>�ޔ0,S���󧇳Ϟ�ᒨ�-��}�!6��Jyv�醊�^_�(�H�(y^����o#����X��3-�k\8�M�T�"`R�DF6ȕ� �,5�;Ҭ C�k���1\������k�t־9�}���� ���QHF��"��t�9 ?��{E_�7��!����](�S��0�q��w�9��=�i]�1�GʦȪc�W�XC�|�$��}q�6����zf(����լml�dz������*�eLD�*�,�m�]ہ6����D�Gw� �g��' A��)�m���b��ӎ���o�6ūvO��=�W�������}��	����z
��z�&�P�K#�^Qץ�_������&�)�ٺ�u#uD�	' �/|�qf�M&P)�tL�x�?�u�����ҽ�����*c"q/�\��YDl2n֢�vtX��Q������ǰ�6K�gVL��ο��Q�������-�˚e��"gb�_� L01�D��ثU�8-��Nw�@�$[�>V,���6�����=����{>G6��v�����φ+Y��	�d�A��b<�)��Gp���k�(�vWu����!5��YB� 5u�8�)7�5��E6��㦚����9x֠"���[����
�֔�I\2��I�Q����dc����c�$$���V���������e�;����Պ�����q,��F�<)_3��i����9[�6��8�  ��؊u����T�]��;���^̠��B[��0�[������ ��c�3:{�a�4����_��	���i���!`x3`��?֞��׊��_���G���!�2(���4��3��Q;�ӣ�H�����_�l]LE����ۛ�Xd� t�4̩/�������Įæ�����s':���yk՚�lP	��񽤒ۨ~�&�Ai2�	�B������yp5�!b�Bw� �9�T�N<�o��������i�<�ț!�"��xOG������dv������a!?����!h����S��b(�#�T���G�qA� �8�������a?��Ly#�N~e�^26�����z��I�A��.�	_ہ�M@��K==��B�	q�%>z�KXR��E�5	�lԻ!ǰ���	5���o����4�������m$����_Y\z`��v���?��Q?X��a_��ׯ�Ҝ�VB����O\��2�|mq���W���/��tk�lҍ���K�\_��u�ww���!9����'_J
@l�np�>Ey�4�a��l��Z����+��y��a�s�!c���i��t��/���G%Ŏ�$�3dY�?�C��I^���;���R�U%K,�r�l�s.����1�F2�����URa֙%�r�Ĥt�x�<�I@)�*�AZ��O!�Ccݬ�h8���1ݼ<�+�G�-���R�:#�#�+N�,����s�ib��W�L��C�<��G�AҔ�����d���������3چ"Wa��
͹�� ���y���j}
@���u���.TD�l���Y?�<���V��e�à��U:�¸�oaΝ,��{$N'� N�w�S������t[A�9=0�3�L��ٱ�ۼdc��UqCiv_�mE�P�o]�wu��͟
��d�	Zn8< |�"P�q.���F���D�0>`2P�p�����7����o�f����@�����������ԁ�F�_Z��SYe���3`c��H�M�K���.dp�1���)�̨��L�[#�\ҳ�5���`�W���m�}l��q2d�C�'�ݨOx)&5�d�H:B���p)�H98gBSdY#8cd5��Eƛph5��ې��Ё�y�.	�f2�{���F�'G1�'�G:,�����4���m��'ζ֜��)-M��i�f�u�ulc�k�-��48
���U�����&46Cr������w�ą��a��%#����H�(�8�|#��{/zp�NsP�����2c�Zxk�d�Խ��qѩf��1��^��I5���
����y�K�#��JUz3e�=��C#�kc�gR�h�i<�;��۾�.��K�%|�݃�,d���GG�7J��s�X�CR}�J�s�$�(�#�$O��(;$��~�Oߏ�Eł�_֤����|���A�N��Q$� �C��'e{IZ�0
ong��'��Ŷb3�t��O��XfT��Y��d���Ѷ�>�y���#��#��2w��MOW���)Nl�gu�3�35�Y2%�=�:�kG�����X7Y���[u����H��_r.���!���<�<GU�����>���θي��ѷN�ܰyi�L�L�) ��@�eۅ1���"�҈zܸ�l�]pB.�:���*ȶGpJ�0ſ����݃|�c�K�����$��a��!.�v� ]��ϸ��~̘� >�#��۔}W@y�i�?�6�V0��"�~���q8�u $g���d)&$��w�bѐO�@r�aWe�]�떿"ӥ޸Q��c��_��n	Oi�:՜]�b��'�:_v�|{���ӄ��Q���8�Kb�}Y� ~�ڡڬ�������Ck�-���k�"���P[����M���8$��H{�w�{$	�2����n5x��1�إ���*V��gt]���"�.*�R��ʥ)�C�ald%@��&�f���qM�V8����ȡ�U�S��F�W ��U֘Rĸ�N9'�l�78�rs�7Op?���<��\>;��)������{��Bܔ.$�hA����ٳM��9�����)? �-�{��eGYM��H�X!(T�΍@�u��>8�DN�{�2�k�υ��JR���������.ؙ��̰��Ƞ[9�m�p_�m+�
:�E�ajHEL���k`��9�	��	�7�H����WzLMD{�-2������٦�����Jw����k����}κK������T�#*����`M���B�;��_��@ �v�����q����|z��*Z��"8��,�o޼H�ؠD��7P�I��'��D9���g�ì��.����#A�<Y�q5��ȸ�[ɑ�,��M�/���?F��ڷ���a�lKF�<I��]��;�[�x�Y< �<$x44����w�o�Jp�"�-�l��p���*Ĉ4�Hy�Q�&�����n�I!��?�oO'�1Ԟb_�޸���V��rcbd���������������J�Ej��Y%��	�l{Yj�Z# j��"i��߇��+�8*C�{�|�	��Vc�4_��pѿ;u\�@�gJ{.���ͫ���d���){�J��l6�Zz�ʐ  aa�J���t��}�"�[�� ��)9�SJ�j�>g�Q���H��踏�}��ک�]�����uŶ� W���A)�$<
|�&�Lb����Bm��E����`xM϶IP���<�`־Ys��68���6��&a��
H/P�պs�n�ȆՔ�+*u�,r;���=�;��hl�Z�5-�@����n���lj��M�g�&��u��}��R�=�����\����u���m��L�1��O�M�B[�^r�X4���kK�η7��;&pQ�I��ꗈr4�t7��G�˼��襾�T�OT��x.����-1/aM9Q��Ay� ��x4�"��&z[}n��D���?����{gLx���l�~�'t9�Lg5�1t�*qB٧�0Ҵ�|�V�0U�F��v�Q�'�\*b�!�*g���ίo�u��H@[kt)�a�������vY���w>��X�W�8i9��A(Kݎi�b�^\o�=��Y�2���C�0�����܋X�"�� �����M�؎:�������fN�6�*:�ܴ�h��Ȗ��}�N����"a�c�X!��f�l��'�ӑy�N]���n���|�$�VvE����@54I�j3sW�O�x��[
�������&H���H�a�X����B�4>rH�����
��Q�L��̘��N��������ۇ��A�D9����x