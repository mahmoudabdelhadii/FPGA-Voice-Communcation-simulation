-- (C) 2001-2016 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
enMN6GsbUv4uB172ptggLmlN4/T+tyQ8yKobOwNov5j37PzSit3dk+OuHOCLnlZKiJ83tShl65Y+
4iHaO0NMyaDGBkjYRcMN8UBQXsUM1d1K5KJOZNsBWucMYMWv1xjgEwE6U3JrZ/7+XqNI9CGUTkMe
yWeQ8rDSf/rtUmsY3BWZxpumMd1j4KsCDS7y4jHwPZbRvzo0lnkT7NH9mijO2AlxOY2SBewzAUG8
2WZAvp4gu2zGn6sf5FZLB774vPy+WyrHOIfQcJVNjMpd0CNCokOsBt8tpt/MZtCEirRmT4ZHYFjM
TdSBeOHUHX+QiPNEszF1VDCXILN7oIqHPffDjA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 2336)
`protect data_block
KejosrDF3lQ0e8D5JBhsKB8dq1rsxvjeYZR3pSF3OM31WsEMrfwlgX6ipsKnOf4O6pR9QZBgLHeR
xeMZ3pCQTpv3nL+5JGu++5RQ7oFJayHACoyh5MDTwGFJDGWoNdA5rAS5YVXV908Av0wHyT4KvvqF
BmL547xhbq2rRb8m786andM4aYhwaWLUF8Hq/T4W55RYma4M+uSk561ihkYIx+PHAHTq06Cs2umz
XKM9XAfj8R2TZWOjYs3RUa1DtOIT0oq0xZEL3Jmsjj/K1TqHMsZxlxrxJJ+QaTVl0jxzXuWx50hQ
YB5Egk+JlRR2amZos5MKtw4WMaRi/H1pgkLrwMeXPJ4O97X1Duf1k4MPCUvC8pwxw7QHbNiisp6s
XbNvmJiVV7kAikAb+vO79rl8VxX2bb4ixS0qh1FWK9keYsRsAnwLF5XomNBZwfKrjVsgik3TaevF
JbnPciRtoScrxKSh6Ur322JDdTimb2w8quFapqwSJLZyqSchaAqywJpHn6a3qhpZMdQH7m6f+CJj
lFNJYEHd2trsxc7lmXZwWeWGm71NnSjc81h+vOwyH5D0I/EP8wpOewlQezVvnB5KPzd8VGrj9q1J
8MXO8QTMO2JbxNHRBm1nTcwgESehO67fAJWfAAt9orwXAR8vTmkOJMrz6E4SrwOSF+jYZKRZ466X
AuGOy4VM8zjiJZdZrBv4S/feJ5qOomrenFLxlR57kK3zgFvnPP0M+o/8haRt2R3ybGcYtSsB2HCN
BeR0tyonVQE6WFEcM3BWWmM2XEQ81CBt4edZWRKFyL3/c+yHpOC8C6HxZLBKmN7vwyHR6ILDOIT/
ABvfcS13cLwGGK+97bFPLLCv+7va0tlBZTqgxWbd4DMXiKQ9KbU6vGzAC3+PrXEMDuom2fvhEhTx
1HdGNNYmEn7FIPXJpyVYAaw7iHiaOsp5sVkGQiQyx/3BVTc1GL+WvIOuheW6e4iGPC1aT+Z0OGCj
9emXyTAvYdbpFOWwcr9mnnQ1DyoSW+ElCdrSIExf7GtUPcKKPoMps2RVRwBpDshP6bhQEBCAJyog
3OpWa6tjAY02XOxIwbcYh+I9LruciSIZioexPzyZA2YtvwcO7SaMRlKR/OdGvID/40Uwzu5yuXs1
mqWAJd5ex3mCm8B7mQ81jPpnqsAPLLbGSr4rjNc3JeTgboQ868ic52nrpXV8scLQKC8jrCgru12O
tfXpaAkFlTYu7ZFtLS2hM3q0ntvy7bRV1s8FmlmRNpcE+P3JrV1OKCEpbrxKor3reWPLZHXbZB+v
21mGrkP5BHkakceL1/ir+VFb+OVufeJYx3Apwth9dol6RGkIfWdIs6XU9tdR4t+PDO9KmXDEt6Wm
P3cmIA+pouKI2rd7iDvHXaMS5mAmu399pohBFHQCUuN1CfZjQ/w9JPien06SFZ5Nwr3WqcwbYuTd
aZ8Tn7Cpg6inC2zQRh6EBJXvTLFlcVZs/e37+5c2WYwhyRbSxg2KxKbHM3b1vektyI3RS7V206fk
SSznPQWlTl0UJyBWUI57Bba+6FfDNlTda+byeKYy7arD7fnjmk0I7urMP0dAe/IRy0ExqCGTQyyw
P2/RRrAKAndXPY/nXQA/PsHTOvvNLylH8jr1xHMAkMxXqHMl61WEh5se1plA4GF50ZzMEAvY24ia
1wF5ed7rya7Mdm57tBDpu9w5tKoe/1jd9pevtfjWzLP0fhGGV1Dsl4BjhhfmMZnOFX7tAAAOTYmW
viUbCdUohV37wkoQNr49lNVokZhHzqDEzaHCN5tUTLM/UMxqI6atcRN4fmS5dEx+cFzNaf4jM1iM
BHKKStHmJs32+FpgJQqg2WyHYfJ50Brk7u94Gahb9QMBQW3BvLREORIxILSX/pm8z24j7GfCo4ea
jTuapfoT1+RtH4BjdWpVm4lpxSVmhHgwa3S/wSWOPVgLYYcq+mUKDqoDI/KZ/hGR2EqfIjYEnM4b
lPymni+SYE9WeqUmXt2Jst7fJ3H/yRaVhjFMhORb4KpzKarVblY5cLllgSe4Il4YSxHjedyXVS8Z
j0YLA2epe13ZdZbjcROqY93Mop368+Cnq74XJ7KHhxkNXW70vNY7ssO6uW8rjKQXPv1OWcngBnC0
6S6weE7qJ0vz9kn84UpKEgYoZv+YpyqJoKybeZpM/hm+BToGRwdcs3jqrOFzCSFOd07JGJZG37LY
dSImNCerXTaOn0B97+5Xf8IuQ0bwF/+9SmQpyE5YFnQLNbfUT6n7cuLBAf/rQrcCLs5WRessy7ef
VxOLDgJ59RnyngjSlpJk7Cksw8WGHPpV77OaO1pGD213Xt9zW0qktVeNGTZVBIoJmVTGBde632Mu
okgTpAx4DXCZFW8oiRM/nH81nsApAUndNHNJXQOgHXQEbA7ox7TDkOsV3Mq0Quy4jeOTs2MIoU1z
4bfn5hnsyD24Gz92ax5X+gQ4UhxaGft+sZh9bFFEeK05+Vi3G1eN35Im5SBoy4OQ7iGyoUGzE2hS
jUZVtJfyFGoSKXwvCi3nDu6737YAZTuBvIn/mVdPXtRK0l4qz5e1BRnyX0iDup0iHP/I4l3J4PNB
ahniYKp657XuDf5V8ctdUHMpNdlz57hDaGkmQlxTK2P6vPO9tEwBRQmMebjsH3mxiRYhqwqK/L09
HLdJflGKmdTr8gyXFaK1FgfvqK6SKT3duZ2wF8ZpEHgRx63SivFPrt8oEFNCCj8TokggVJuhwpqh
x51u9V6kUYUubndukyrco/HQRbcoAqAZiikNB4lYLcyUHxUu0PaNUas86JDLbP7UPBzfmcNh5xcq
3eM2CcZzFcaRIeB5vsquWb0YI+l2O2ys1fhDf9G1W/dq/Jg6rUDoTKWnt59mzQOMx75yClFm7r4Z
cXpmjbmiCAWjFkn03zi3wWKJ6j3w3zOhSQVE4sNcYDoG2IFzwfzAxNNw4sW4zxWGfSy7SD9AoDZl
Ebat0tMT0IducgRUibCXm+yt0AnDWkCSWO4TlKK2ppviiQyXFBRjCIkHzITBWiwZDOKpFCp+dIPh
RBuXa91gCfboJv6QP+rlkIr8P8S6RnFR71UsJMGW6IAXOVWpt/uffuAhsz7HOr6qTc/49tViXDE=
`protect end_protected
