��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����N~@#�k�0!����+��=L���0�ԴZ�2�Mc���ZO�����=�����վ�	"cqw��a��TS[��{=:�����K��-�մ�(��k��N�-� 偙O��QZ��~rL'�x[�i,mׇp���O�I43��4d�,�H�����SN��d���3���r��m���̨T�I;uj2Y� Er�*p�Q$Gm���p�V�`�2^���,hz�<p��l�Bxt�5��s��\yq���#�@W���f:m��T�	,*�񞭋����_��㧋l�	�\�:��uGd��PǷ��N�I��_����Tuv� ���us�(H�~�{2H�:Zor�Q	#%�3ˠ!��iS��95�,?�.���/�F�i{#���Tp5����Ҥ0{%���2vpn���X�����@l����3dc�ק�3	�Ed&3�ZN O���z��s�yxӡt��v*}ԫy nj#��lc��m戭k[��5)�A#�����8�!�]�Z�s�M���t��w�!��'ÒE�rv��Ϝ�c@<U��\tq+��&|�&X1)C�����r�A~��B�&�����s�:n{p��͠R�X⺂L^��R����c���f��J^?��ܣR�O 1�rV���:��T�4���AD����˩�F�w��)Dm�O�b,�a���1$��c��7t[i2>�ޔ0,S���󧇳Ϟ�ᒨ�-��}�!6��Jyv�醊�^_�(�H�(y^����o#����X��3-�k\8�M�T�"`R�DF6ȕ� �,5�;Ҭ C�k���1\������k�t־9�}���� ���QHF��"��t�9 ?��{E_�7��!����](�S��0�q��w�9��=�i]�1�GʦȪc�W�XC�|�$��}q�6����zf(����լml�dz������*�eLD�*�,�m�]ہ6����D�Gw� �g��' A���FX��\өܹ&�6�h�Ð�$�(+��埧��= Eza ��찠pr[�c&��nP��x�2�TK�M�V���3Y4vIR\������ɭ�1՟?4�_y�y+����ƄJMm����@����m�����c�t�����:ud�Q�����T4���QxBŎ��\o���t�*Z�$�*7<�t~eP/`lfhg��6��[nn��#<����n�D:� ����4��y��I�I$�c�	ꈞ����G�l�\a��~�a-�]EA��|I�{��#�N�e�R�+Ø��fyz���%]��?��*��XGa{��!�N�\�$� �˨T9,B�-��Bt�S�Ft4�V�8n\)�Gc�B�b��5��]Y7�1��ȴ�OvG��Κ��ئ>�'�_��M����0��*?���$���aο�Ԙ��	e7!�
������3�>L�zcA���ฉQ�!8@�3nd�~����PU �`���1:�hr����+��S�w���"&�(��B/$��]T�ҢY)x�+��+��9eC!?�%)31�Q4����
@��� ��pz{%Q�$��ǿF���0~S�`L���;�����8W��u��:���#!4b�hn��JBl�	� ����:ӊ#�v��p7}`<��-���U�;���3���g���sG��-7Ԧ~�8���$;�X��&�}8|H=H
�O��X��W���b�mh�!���p�7����J�
�h��^Ly���Q+����?Z�2�jh��B��$��\�9+��|f+�f4��+�m;��×�o�����Xx �	�ۆ�,�ct���K~�"���Ob�P�~�B}8�*���{�Glj>
�c��[&�&���XV�#���}7;1�%�}�F�>O.	(��4y��d*9<���m�W�v�ō�ʱ�wj�W����=H1C{���4E�Q#�UB%ѣo��Q�rD���z�0@Ԇ�׎L	��	~�*���i��K6P��#I%��kD�d]��b�[��	j��k9����j�(uB���YX}v9}�18�l�k�Xg���(U����ϡ<->�%oe֖�L�!���H��`6]�Oc�yo$ ��`��y���癷��y�[ɟ��O�s6��h@�T�5]4�-�GS��$�b�Ě�����zY`��.MI��墟�H�d���� �(M�_�`�c�����>:n����@��V���-����a���Թ*��eQ6K�Ÿ��o�=��x}l'j��#�T$���lm߭V���8��z?`�I������q^	C]Z~YRvB�]b����L<v�U�n�y6\^*] _�-�I��.�qm)9Jt��Rk&��t�|���IY�U�˶I�y)XA�n7��I�5��D�u��$IL��|���&�R'bd��g�*qf=y�i����r������m���\o�S����Ռ@�us�^�{u�b���ޱZ�@�񋳽
	N\��t����B�i]���`)"Vyks#(�^b��ބ���1����qP�TF���{�ȓ6dQ�Z��Q���ײ�&Y'�-� 6:G�s����\m@㽥u�?��rՄC�m�����4�쮪����n����>�(4]�8>�|�[���H�h.�s��BD��]J��芴��%�.ͳoX����~�`��i�Xݠ���;�%� 5:��q-J�%�x~�͚�h���3�A��l��w{q�a�������i]���`
��Kr�r�I����Jsr�G«t�
a�=2&�����_��@^Q��>ƳD:���cq��I�� ȧ���ր��s@2��TGO�#��y��O� �9�'
��\��������}$����z-���p���@y�d8o��Vp�4���HBz�1G��%��1jh�ꮕga�2��7���-�#��Ҽ��wq�-�뚲@���`�^�/�@,�~�@�>L}S�*H�GO�����n~��\h�ňW�o7W(�Kl)���-��nϹ܁3�0.(��C:o��_Y� �hlF���|G�fW@��#�=�w����0i�A)J黙$�V36B���N�( ��93��0�?0�ǩ*�<z�X����Y�6�皊۠�U��c9�)�;��;���~w�y�W�i#�d�Y��O���[W���$B���I��Ց�μ�2���&��G>@*��J+ě��1?Ks�M�|
vg˩�B��Q�\'�'��ñ�����d�c< ��A�e��P�cqI���7(+�T�@>�!IM{I�H5�aM�l�a�N�\�2�q�j�v{�vC��cJ��PD`�`�f�8=�[�����O��E����&��-�aE[�3��~v�Н f6�o!F���<�%� �J5Od�Zsu*���1�