��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��,�y�}�ǰ�=4d�H���`I"��W�`r���T:tB�T4D�m�)�	1��I�t��
��8(�8t>s)ו�."[�漆���]�~�]��;�O(1#5�-� 偙O��QZ��~rL'�x[�i,mׇp���O�I43��4d�,�H�����SN��d���3���r��m���̨T�I;uj2Y� Er�*p�Q$Gm���p�V�`�2^���,hz�<p��l�Bxt�5��s��\yq���#�@W���f:m��T�	,*�񞭋����_��㧋l�	�\�:��uGd��PǷ��N�I��_����Tuv� ���us�(H�~�{2H�:Zor�Q	#%�3ˠ!��iS��95�,?�.���/�F�i{#���Tp5����Ҥ0{%���2vpn���X�����@l����3dc�ק�3	�Ed&3�ZN O���z��s�yxӡt��v*}ԫy nj#��lc��m戭k[��5)�A#�����8�!�]�Z�s�M���t��w�!��'ÒE�rv��Ϝ�c@<U��\tq+��&|�&X1)C�����r�A~��B�&�����s�:n{p��͠R�X⺂L^��R����c���f��J^?��ܣR�O 1�rV���:��T�4���AD����˩�F�w��)Dm�O�b,�a���1$��c��7t[i2>�ޔ0,S���󧇳Ϟ�ᒨ�-��}�!6��Jyv�醊�^_�(�H�(y^����o#����X��3-�k\8�M�T�"`R�DF6ȕ� �,5�;Ҭ C�k���1\������k�t־9�}���� ���QHF��"��t�9 ?��{E_�7��!����](�S��0�q��w�9��=�i]�1�GʦȪc�W�XC�|�$��}q�6����zf(����լml�dz������*�eLD�*�,�m�]ہ6����D�Gw� �g��' A��)�m���b��ӎ���o�6ūvO��=�W�������}��	����z
��z�&�P�K#�^Qץ�_������&�)�ٺ���/��U���WX�wK³��4�d{B9/��&�	�d �Y ����6��-�X��o0O6K�-آ6�F�,H+B�*�5	��~��6�q�?T8F��Ýt��_Kf��b�Myz}���%�l���)�|��za�ӗ*���>Tk��EU�[��2�Lu�uU��=��L��Vn����$a�9�f~U=w��h�l��r�7eg�1���$��=?	)�Q��^��(�OɦǤѲu����u�r\QD��q���ts%��2��_\F�H��,��gm��1��&^8��,��������C4��xi���%?ܡq�q�(R�N�ff�E�\,�t]�2rđ �J��$�i+�7���a�"4���v���\���LFsy��,���i͆)�@Z��N2YA4q��a�����J�](�6x[9T�����u[��E�Rj�{%�O�|�Y�S]�����GE�O���#<C��z�<D˓��=�e�ﻳT�<��)t-Q ����_P]��M�#��5�r�`q�����i~�������P�$`��v��"K�����E�!?����2d�V�BiFAq��a��o�J���9�]p��D+��P�x�&�*D�r�Y�AEa./X8�j>�O���:��X-RXn7�]kNҠ�q�՛���C5<}�˱�]yY`�u�$�"r��7�(� ���c�}5��>��L�dX��B��¹��b��>�������>�w4V{������iϪ�~��3�E�MOaq>.
|aX�W@�� ��!UM���#�Ej1����zX�ѫ8Tʠ�u�-3R���}j$l��R2��"˓Kf�u�C+T�D&�w�j�l�W�0\*3�	�Y�v�����C��-�D^m��T��r3Yf�v8�(p��йL��ī%[�r�%��מ�(@�����#���;Z&�|,�]T�ҫ���Ӑ�(�Q��"u��;�׺�O,-I��jr`��q`��O��*,�x�#�t���e#�SyM���@�湯��'�D�9�V�����f��-��ġ��o���+�����Z7�$	,���)� ?��l��tj?�d�l��G��/�g���oH�rU������}� xu�e�>9��s�M���#-�����B:��� �������S2�P�[)�Aj��|�ͻ>7w�������W0��R��u����1�h[8k�S�Lf����*5b:�2���S3c==����3]���\7U�i�ŭͺ�X��_�vU��c�"&Ų%?��+�fx�,zn�8��O�2�k�ky�o��{)�=�bUL{�>�%yWDt��O�A{�|l�W}��x�Y����+/�шրWW�4k=%�u�����˿��줥��awj R��z�����g����;��:�<��R�π����g"oq���y�K�ie"\���4�?�L�'"���I��
H߳b��D����s�0B�Ԋ��E�Q!{įu�U��0��V��ĩEDտ!o�"{=�ۀ����Xu�2�wA9<�dQ����L\��	kd�������痳!����D��/�4�*Þ��ۮ�����Ó`,~����7�,�{gӃ��I�J^TЮ_�3%��C�U>R�������"\Uk����c���v{��j�#PC�J\pZ=�QO(�9�Ǐb�㩷\G��q}��ƾ���:��ߩ8��I>y�E~y�]ᄈ��Z���ȓƎ��Mױꍇ����C��Th򳠝�7a�ԕ��.�!�D)#��)Jed���;Z��i�ۂ�;?�nύӐ��5 ]�Ƭ_�{@j��@\-zMg�T�=��v�y5���mH���y(�X(?+�s���r��+�@!9{kw�N���0������.�K�wp7��qo����C�C�g��;��Cv�N�V�
޿3�´�­�}�X�������N������]ͤ^���ALT"�CN݁�Do;�i����~j�ãd��/��YX����5A"�hvt���oHI�J�M.'�Bƽ^��!�#P�Q��S�t_��=����f��23R�=[P_�+���Z����10��t�(���p���Wx�`{�e*� \�P<Ku�>���E��U���w_���Py7"H��r�[��=�I�c(`sN>��z�d��{��z�n��dX�٘azg@��wL|$�Ee�W���s�n�	zU?�v��A�䑡FJ� �1����TQ�o��;_���:'�
��i����	�����V��ut,JQy�v���m�z���ԋ/���y;�h�kſ�����*�|O���r�z��h�y�<(`+ᣃUSe��2�f��9�6�I�ۏB����K՟rL� �����ee��7��~�~��ԁ��}�w��2V��B�PY�P�\(���E՝��{s��hd�N݀��Ŭ���p':�/`��M�ΫF9���B/X�al�ȱO2�%��f����/Z�������~A����{w/Q�v�|)���������\��@0�o�Y���e^��cU$G��1&���SM~�1��	��#���i�S=�4Y����#c����C4{�T�A�:L}GؓZ鑵����'�#�?O�ܵ$�C�!�N�5hv�s�Ւ3��|�V��nN�V�w��&u�M�	���k�ܽ�b
�54���b< �x�p�?�_���)��ԏnG���nU����)������پTov�׻ZOs�V��V��!e�T�����
TI�}^ve1&��f$�oם5�SY�O=Z�_ω�����(	W�X���O�Pޢܦ@�K��:ı2w�2���l�s��6��m�*�1�֩8��_��c�v��㐤�rW5�@����m���J�m��w}��t������9�Sg�9+Z<�'!V8�w��)棂?�cͼ�gq��� ��J�\e�UJ��;~R%���y�cP.<��<6X�h�24�"Ӭ�U�2�����
X�F5�'��uP�T���v�BJ%y9h����Fjh<Ӥ�9�V{Z�9�r�rx���W1w���F��F��n;d�c�_[մZB?�Mj[AC{��鶐Bt^g��S�����O��)���ZԢuB�����k�7���0�� N����@�A>˧ux�f"����S�P�2�y�l�7L�+x�>�%��k�����Q��}j�y�"UuBݯ����F<h�z�O�.�Z��� ��Dqn�#5<���iz��ɽs+F��B��|�xϨUy
.�}�$�B%�[�_C�%�x۳��h�i:\
p?���ǣt�ݫ���$��b<Ac5Q�4a8�#�l�΄t�	z����(r� �FVChMI�I�xOUl���8I��D��o"�)�D��J,�0}:���_ �߾S�@?Q5h���LŒ6\��Ԩ���2�~T������	����\>�S���T$�K�1��I��[�5C�D�@�$��|��{�b#Q��E=�{��ݠF�#A20q�rF9��*0�R"�i���K�̒�ܘB�����Ҧ��߹�a�02A(ZA4[���1�cD��;�g����<�vc��%!e�� +�������K�QO0ˬa��a���=���ѡ0@�:��_AYN�R�Z��m@m8K9�^lX�������M�s36��4n\�i&����z��%���m�^�@��OA�Ue���#�tT%=K��NI�����x:`�ʦ(����H}����������������/1���cez�Z�0m��L��3�+�����6s�~��q*_R@��"CJ��k!�_�Jܦ���4
*�X������uN�>7q�de�ِ^�����qWnØ��VQ� �-G�1A"���s:)Q��Ьj�i�#�>�Ӝ#h�"&x�>���4��x�������ٵ�f�CYz^���悺[|be�:��6m%�%�Vgv�����Ȫ��T����m����+^X����oخ{m*�'4O
j�VJ&�n�.-B$�ڪW^��䜖���1��75��6ʪ��g>�f���]�㥫��nx�,�e6���ٴg.|�?p_���طF(�q�i�^t���JZ��K�+v��d�M/;F�/�ܞia�t�Ğ��>M>_�|��8�����vů�־�,�v�Ϩ�����E&6�P�˼�TTa�LI�\$�����%w����+�\�q��$6� �kp�\`7=
��0/�Ƌ(}�ȣ����b���K��G�ںI@4^��@m1���VЧbR׳�SK2�V�}�m��N[����V�ku��nVUm�WzBܖϓ��?T���������nm�i���&����Ў(�b �9��yt�w�t2�1ak��][�u�w�P���c���߈0���#	ꛎf|}��|65ݽ���KWr��פA,kg�
 %�P88"�d`�����L���a�I�݊9!�6!��0t7p��/��!E��"��J=Y�#uR.}�E��i"���.@
F�L�ڗ�ax��GbA�П����-[�YI�U���"G��@R�CT�˔҇�*��lG$�B����*|)7�.3��lғ��!m|h+��:��C��U��f�'��U�(Y���6A��(hw���8Z���_C�5�-T��ВQ�I�x\Ab
ʅ!��t�S��&�����K!6@ʹ�a�S)�n��t5�!/YKn/�D%��åaΛeJ������a�m<WK���Ć�I�gऐ�/6��)٥$=	��)��ӫ�_���T��Y�)Z�82���`��+����+9���.�%�༔���~+9I?,s\���RdƜ]AK������o4r~�����Q��S�;x:�A%B�Vi(	H�w�}��0�E�J�5i9��R��mQ������ɽ�Ts�WA]�L-6M�dٕ`4��q\�`|d������ԟCɥ?t���Gq��9�xR�����ѩYD�3���ѡH�{,���(1��A�E����W\c3'X��k�A���\p�~���@Ӎ�"c���K^&��b�b|�Zp����N���	ʿ掷p0�=����<�D�}XW�W̫L�D�;!��wpP�%8NG ����2[t#�+�����[yx�k8��w{��E
��c�2�(L�߆�r��e*h���`ȳ��I�av� 7�0{_���?�,(#K�~�J�s�0���f޸�T��By�m�/�$�����F[.G�,N�*�5�wxu�-i�1y<nQ�x�7�U(1-����/���"�M��������A�lz@.8��e%{ؼ���*e�9�m�$��}VF ���rq\�A��{�M�r� ���r���>�'9_��5$��G�z��!��o��:��A�G7�m�p}�!���F��r��0�w�`�]s�1��_G�#�Ћ���	c��?���}J{����@��պv\BT-�F���j ���Cd�P�Kvqk�8S���j�oP6��2%[̝l��I��+ ��0�U��_�y�w�7I5W1�ҥ
��q���46���V5�߆B0f���ǃ��,z�r��3=�L�d���]<Vp�T�$�M���Z�F� *P����k���I>D
�[�}�n����{�pj񠘐��>��������z���5�ZK�8f�u������хy�� �������rd�P�,�P����Up�ʻ2�iP�M���H���ߦm��׺��n�t�h7�j�#7%��Efh>�A�^�m����(�\Z���� Ӷp5vS�:Z6��;�t�0�g$���*u)�K�'گ����aY�U(7b�J\����yb��	��oˋ�8RTY�,�<��s%H��o�5t�Ąn����r�7
��l�_�D��'4�"�S
LS�V� �-�hOzv��Y�]�"�s�����r���]R�"A3]7�`�~;+HyF}��*d�V�y�Br��(�Y{ׂ�3��E�Ţ�L���Vz%� �@����"F���s�#$��m�c�Y	���[��
�]�����GmTVAK2�3=�Oe��z�a�T����\'C�:�>��ߪ~�-�x���Ń~��=�ܲw��\bu�dIF�=&����C̛����C<ջ0W�s��]��Jb���c�ۙs�A�	9w��b�Sa�4����m��B~"C��h��>v�O�}q_yN2��.p���0怀O�.$n<�tG��zq`>��~��)�� �q�6��>�!�χI,�J�刌�C��_D�D�<�o= ak4kt`@WҾ���EQ0�U1��%�q}���?�2�a�~Qϡf�{�-E�ufl��1A]��_ͯ��p�Pt�[��5m��n><����Q-.�CJu�b`��0^BJ�M��D�e���cB�]c�?S�L8��p����ch�S%3��Y@Lƻ�(z�QD,��6[Y�ъM������}�qh���)�PrZh�H��:�I,��g~���%x�٤<+s��z?�^n�&х%��ȩ�@o]�X��n9�4v�^��K�.��?���R'�!�UC�s!2�[��Sgg����䞋Q �C���(\���`(p��p�A��E�Ӳw\i�}B��+�tmK���������7�#��/oLK�q01:���]JͰ��M��-��e�T��2�h��n�;o�z�D�C�D˼���?�* �ϝW����(�rP�3�~���l�.���)ۘ��3����l�ܛ���*z�|dns#HHN���[�܂h#D�,M(3e��)sK��rs+�.P�"�J���a	*.]������+��Ԃa��/�lz�<��p��+�w�����@��~L�&��jTl^j��0�TYoe�&�yTnD���rl�����'�B�@�8�OJ�8sp̢s1)��д�ʁi9�����O����:���:�B�>/����2����#z!F�k��||��XW�I!Z�0�N�� {�Ǝ��ؔEa!��n�}���$�*e>�TR�<�d5c.�r�����J��w"�cx#Is-�_�"ٝX� ��]�)�ΐ������?�l��w��֗a���[��ӧ�ᑜ�i� [ �q\���A�' �V�'�w�u�8%��%��;��ǧ�ٯ��XB�P�)����L���YX���� �kO����]�Ǩ��ctN�[}��ӣ��+�wv"M���~u�Y��a5�g��E#��W��ژ�M@`=vQ���q�	K�p��_�`�����A/]k�$���Ճ��g}�ZS�KX�>f�����۶�o=q�v��RT�8��d=0��ڷj0��u�Ƥ/��������Ϟ@�:J����?��Ƶ��^���l�Z�R��D���Çh��׫d/�q��h����^�]���E��C	���㒔^?O�^�5I.�e�9%�%t�[T�Ɖb1�jt�e�s�N�,ѳ[?O���S��į��h��vͽPɗ�Ly���=���j?�XqNK��:Zn]s$�Yz`���ƻ'��"�̛h~Ǖ�0�1��ڠ\��7"�v2�;*����e�QJ� �V�s[�Eg�o�.�`��1���pq!��@����[J5A�|t*�&��,I�^��&t�%��$O��Ha�6W��XՙΆ}��t�j�K�ո������1�Ϟ��4T1C�4��'շz����x׈����7aL=��9�B9��ճ͌��K-�C�Rk��t��x֝��i����2��4�@���jr���P�����Ki��I��{Uz��<�_�04w����mcn"��=5���)CU0�}�-���i���L�i��	-ŉJ��3�9A�yY�p0��OX�������1D�D�y`�vNK���Ş�����t9|'���I
��\w!W��\w!���98ݤ|{$�B��-/Z��!D=&ꇎ"���Mlu��^w ��z���P��?� ы�����n_jҥ�Nԍ�z/����QJ)��5rժ�w48:E�J8<�Z<倜�u���>���&a�j�$M��v��Ќ�
h�Xl�i���m�Y�&~��&��7���ث���[�?D�0�Ikr?���^�2Eg��
���q5S iD������k�ߧ�ݍ[��T���9��0`��(^�\g�-a�vU�|�k�8�K��%r�{}I�HK��j���k��	�3�?Y�ŕ��aNԪ9���{	�����bN�K�[V��|=Z��w��ŢlI�'�\�H��~�S�����2�M{����S� ��[s@3p�؁bJ�]�T��h�!	.���|<~�e��
�M�+��?=�֙ā�2u�ԛ�C�ic����.�S�V'�Q�ri�2Ud�A�хI�N�%����R����a5��)�@1��D[%Aw�l�vW�g�s�U�u�_�q;yܓqJ��^N��6*� _����� F�{/*�pZ�WĻ�
��D�����w��FٲR��`ul�K >J��/<�GV��Rꦎ�l�4͝�S�{ͱ�6�b�f���ݍ��C����˜҅���$�ҳ0I�0�u�X����*���9?���-�RO����2!S���$�7`(��6��J�ŁQϕ�ø��d�;{�۔��aa�|Uy烎��?/����:u��Ud���_�n�	����ZE�.[f�b����e��BO���/a��ǀ�@��1(;lb�������#2hq�o�������%|���/(�	*=�ON)�dUF�����)[�.�	��yo�C�婚*a��rV�#�p���2�L�1�g[���a���J�D(�&�*��ͺr�Mgv���4#���Ă�9~�VmȂ�&��$[��?QV�>��Iɮ�|����3TKP9~��4b]�:i��ڞ[�i4z�϶��,�w>";~���?'���|�Gj)7����	)�e�.����V���l!e��Q�0���p�"v�7ge�"n7�g><=�T��� ���x>�d]��Y�^	��t��ƝS,z<� �#�����f�f�Cb$�'f0>�����f�4|O�e��X�:^�~K���� =D�U���A�)����U�1��
1sNkaH(��ǐ}��~��B�汃Bo\�[�)�Q�����!97�����dэ��7��s1<�q��$����=�'}�n����;N�y��������5�g����:���U{�7�T50�Py�
��7���h ���p���C�b%�p�PF�4hT*B+�֎Q�l��1�']�ώ1��^��
���q���}A�B�R`�vm��,�
d�NF�q�~��B	(���(�R�і�� ��1>���'/J��`���-P��3�@� 潈'��f$ �3���.pd�]~؏��
T�O}��_�\H�N{�bAh���d�a'���F�O��'F_���Ptu�<����&Qe]��i��vg����@Ґ�j�i�P�m�Na=+RO��g�P�����rX�G6[��P�i�������7��ZC˭U� �F�4��џ&��"�I:�E$(����w�Z�kDb���-@�����(�	�.�P�j@��P[�Iާ'����JA[	R��� ���e+�������v'���T[fǹ%1�6v4��5��T*$�"�fMHq�4�=���+.�lQ� �@��M��7��@q��������F/���$�F�κv�8u���T(ǀ뗹���[�s!��
�&�A�-��s�2R�y�VS�Zy<8z�DS%SM�c�c�c�,����ՠ49a\��$��j�X�7Jq,Ct�H.&_��A��_ѼֻA����%:dc�Al������1�S�s*��ڥ���v��CPغ�˔-��j����ʥ����b24D�"�7��P�5��z�̠������mZ�n��Gі�ݧ�v���^�Xn�pB��W �?ߘ��qD!N���8R�5|I�/^C��t�p�T�_�	<�|�ƅ�rJC_�N�D�@B�cß�!Z���5H�iyo3�]_��H��|���""�V���4~k��һ⇉|� ~�����6�L�z5%�͙��u��q�D��W�9� It�W[b��{�{���1R!�
����2_j��G:��Ti�y=������YPŜ?Z�*nhm7�@���
�k��m��K��x��y��$�Vr�Ї���1pa|/��
�c���!U���=snx�`�|G(������Խ����V��T���Wt���i 6���k�o�?�B�����ܥl|�]}
�ɂ����O�j�	�EIgsn)4j��&��ßl��M�!�S;I6'��,����40s���O���6�c)��4���ⷚ"�,�þ#B>3UN�W���v( ����Ю�gH��Y��C�^����)1����� 4;ݣ��l�e�l�2�^� am	~[�c��k\��b}���}%�b*Bs�-�j����w� � �^�Bw��r�/�~�*�z�g"�� m(��f}�*����ͽ��uG��,� �5�x����Lɥ��\���+�E�fK�������_2�R��n�@Tu�^�����b`��-y
�jIBɱh�����&��z4��g][�p(�����7��/�Z̴KR׺'�[���\gր�-ث��dN�*���.�d��bZ�?ҕ�W��uH,R׸7��㕃��Ŝ��r5��>�M��q��� ��ò��%�~A��4�q���`�L�ɼ�:|<'~�ږ�2S#��c��?b�gPl�w�rG��F2��}Y�KF�1@�{Ҁ�&.*�Q����{�/��NI�TɊ�.%B"��箏[GGz���:�1�Ay[��>~C`�,��R�&�]��uuf1�A�� 	uf�~�Ѵ����@�̢T����<8(��+�Sd�>��cɗ�1�F�a�񒿂h4�Mw q���� F�����:f�� ��Ƨ��T�q���ؿ�(�'��">r���!����������lu�LV�|M>g�
S��?�X�JPv#0���^�LO�u۬�u�(�J��f�J�
�A�����Zk���f̄���6�Rk0�0!�T������]�1��+\"�J���P�aO�=vХb��&�1� Q����]~9Tu�n���I_ps~M܊H��$D��
'�N���K;�䓜�j����]�
��&?�,|�Lq��9E�m�g�{�Ē�ᚸ�.�K���ri��JW@,XERҠbt�D-�:��8��&�aY�^F��5�`��3�� 0�<�5�i����B��?�Gȋ�����e�V�9pF❡/��6b3^��b��R\�&k|�����hۨЎ�����mf_��V�:n�#
-��M%d������(��&-��m��P���Jhu���ߜ��E�?�n5���M^W�0�Tݠ��p[��u)s�8e��r�N�3�ȩ�_���5�����4�"���	����2��~�<"��[��4�R"MI�S86�ȩ�� �c�d�ѹ���Q�"{>�a
�se�\���@ړԦ�G
�,�Q��|��נ=�;O�����q�}U�������H	E}�<҃��d̅�g�����E�>�������{�1���P�b� ��V�=U*߽�!q]��IC+���Z���oH1X#*m��E�k�ƕ����vjD��W�h��=��B�����iR|�fհ!.U<��ڻ��gm
.�Z��n�9f{q�E;�5��EQ�y���h@�`�l@���;!c���#������E�o/c	ث?��L�2�U'��\l����X�ǉ��hQ[6�l��$�d�F����÷�G��P:�&�m�
�^�ǳ��^�;��B����|i�-ta��د�|m�jPTWX�X��eO��d��Q+��e!�8������S2�A�?��C.Ãx��f�A����BR�$���Ǿ�$�AZ�|����=��gf؃�7�+2r�Dk���t�ߌ
�qL��5O���벒8�O�(��z��%-f�ּM�	��A��|�8jG�
�~I^�^���`_��?4�GLM[���[�B��^���gȈ���Nw�h�K�$����N9,��8���PWL�E�(FvH֦�jM2c:Ⲙr'�z��p������A�[|�����b��`R�ǚRZƀ�d#�b���ظ 󻣻�a�~�ߔ��C����uA��$��YHG�D��&���̱��:��.fh���TB����C�O��,�Ȇ=Lz���>釅�o"������KaMd�ֈ����Gf,��9N%�ᨅ��	l���V%|תWuӎ���YJ�����;n������/1�죚L8��E���2~�=��!	ŵH�y2�c�o������Y���*W�HG<6����[�M�~_�y5g|'�0eƞ�e��d����3�2�sAڜ�}�+����0j<
�������+�5�n�l��k�l�'X��y��٫��e�!�Z�@���]�rAt ����ޭ�����XT�A��=�6���8>�BM0-�b��R��R�Y�,!���Ƈ!D��	�g�WjW+��ْ$.���TRw1�ֱ������)��)$�`�ˀ�����Ug�sP\\>o�,$-�c��Y?�3��Q!� '�N!���Q�3t�:�a�������R����锣���ȏ"S�+����)[{�:�7ZmB{���yю�~�l?�۱�^C�����.w]�g�(Y��)ҥ�Q/�8�����@K���Z��� 6�Y���R	rQ���������H��-!<�MJ˝�M1��A���ڏ�ۊg�j�Wҡ�/��V�BB� |$��W�7"�0Z4f �q~��i>Qm��̯D�D���0�(Ģ�أf��#�b\����3�
0ȧm�	g��6�+��ԓ�ἲ�*p��=�剗�F�O���
T�"��\�:~ ��,g�Ȱ������0�C���'�;���H;�LzF�D��C��V�[�i�O�P�g*�k��N�
��6㡶��V�t:O[叕:��?j��.q#R"�3�T��u
����@T>�[����?(�]���QGla�) ���[��(Ɯ]�c��E��IdG��r�$��%qN��n�8sɏ�9!־>�������e�I���FHx�� t���a��)�6��;�b��D�)�?h.h}��� }Z�x��绝�İ�/���)X�3im���]��d����v���T��Nb�4v����W�ց���},�l[�mU�T�OAj��ISğ���t�%8;wc�铊U�����5[��҄��	�-�c>���Uv4�X��3
�[ ]�T[���Cm8�h��l0A���g,l	 \������tGz^$�'�����G��k�*h��o��3����Bp��AA��.<���̠Tt�x@���'�T'f�j*i~+ P�F�������^ʶ��������. �Uh����>�w(3�K�Ѩ��J\jKWN0�{/
��:m�y�ɧ�MA�-��m	E]��I�-_����m�7�Es�K�n�:V�l�ǜp�T1b�?�jeRA1�Q#��s$K9���k8�����`'�P�벢y�Q�JF|��>�<E�;��:��+>$���ľ쥱PGFgV�Kt���/�I�_Z����Y(��zK��_�>T"q��^��
��I��N�ˬF��=�b��K��f<)�\�G�	���/�}�	�x�v��J�0�"��j}�q���Xg��i*�H��A�i.-	m=�E���:ֆr�1*��L�z}�IgK�O"|�,��(}�Q��搲ߏ���|c�^�'sj"��� �:������.����Es#�{��q;� w�9
Q�4ƕ�xg7�t�1��0�p;J�ⲳv�8Wk�C��u�1�kr'��,o��^�qS�䃞.s�?f�O� �H�K�C�����)�����%\�m�{	~J�Qh$���g�)C9)��e��DV֌�ڵ��pO�L�>*�w�Wp�o�������Q�n�g�B��� ���=�%�w��;3\k{~BO�D���B���Z[����L����
Åk�C�QT�t�GۺYJpٵ�E]�G��'�M���K�6qt��)��Jy���)�d}#��}k�������\��y;���!�|U��$��CØ��}��AL��uaH>��:)��Y�Hl�f���-|/��7ph�����&�X�?���)@�A"'-j1_:j�
x �9�g+_�(9����1��x7��<��$[D8.-��<Fk(*��D��kP�;D����.��V��wˉni��1���p�L~Dw��g�� ��46���l��$�f�#F�`yn]~kC竵+���+�e�U�fxk�2��ʆ�^
���� �Z;���D��������epiOZ�m°x�-	ܩB'x��đ����l4�w�w�PO�iJWJ��Xn�Ӄ��+��u f�z��/�i)!"�j��gm<�:������L��܌Iцxv�_���Z���O�w]����y[�@�����K�2���	�\��wUug��7�{����@T�
&KB�z�:���a5>�-Uޏy[u�R�{�C�ep��̻|]��>�~�t�R"a�A��=����17���V^���ߝ�e~�n*bݢ�v�Nf}P_��D:4��h�Z��_������ ����$˿n�6��� ��M�V�뤺��8�u$zh�K�����kBƷ�?_�_��$��Q�i��}j�n4;�����b�DAt�i);	��DzJ4��Z��v.�J�0dV�h����|?�x�*Z�x`���N㰣��#�S��a�|��!К&_8�[��%�ѩ��F��Y��"��:���h=Y����ao�*�R�_��Y��2��@bd��9$�hW���S�g ֵ|_e�1K�/��S�8��X$ʣwu$�
qu��S���� ��S;�a�g	 2��y�#ط�&��r���'�%Tu�	��\#����[���7ɑB���mԄ6˿)WW��^�I��X�菝W�[]��l�O��ע=�q��G�-�Yi�Di86�#�05�I'E��ɉ�s�bpC�Ҕ��fP/0󽘩Kc_�lQ)�_�k�*Z*#�;'�tT|@���mo����!֑����z�p���AI�1�\���%b�A���$(n�Y令�i� ���.��KK.�����ϾP]I����@ �axI�x?��#g����-�ǪӒ��62aO��ш�ɀn\�~l�(�F�D���e��R��{6²�"d�>5C]9r�.�_'*R�$�*�6}�Oۑ*����Z��f��[���$dA����p��Q�K�9�C��Fc�fb�$��VM�d�vÊ��D	e��˞h�'m,c�ag5�EW���������Ωi^����MXU~�����]��2�ؼ -&4��_n���!l�/E�XQ}��]�v�,�-��a�Fn�%�AB&o�Q�-�j�3��'�z(��hײ��ܻg��!m�a�n^(%�̙��l�͋�����,5��H?+^0Yh��gJ?��#Q�q��/BB�	�p�L��\�[t�]�"�e,F��H�׾"�����J�v�� N C�M�y�[?ؙеI�����*!'�P}���H e�!�BS|wE�hl������9��f�rw��8.�G֮��QԔ��"�pq���a��-Zs������S	��sI�ה!RD$<0z��T#~�޷ųP3���L�J�� e$Ղ,W�*�A�9���h��4��l2Qw��F���B�M3+�i���O�Wi�<��/�"|i�N�}';�3��`��\�c�F���M�7�~`y8껑4��	CǓ)%i�c�G>�M��:h��2�d��/�f�����jg�,,�;w�&c��+��}˄��o�@T�	t{�}P�ĳM&����A�}��I�6�R�Z]*)= ��*փ��V�d�P��9�Q�Z��v\A���>lm�V�����7Z'&�,��П'����p��\�9Wk��Q���?�$ĵVu}�۬����=N︅� ���[��-�(O�G���9��L� tl٣�)Q����va�e��@�יÅ4�5 J�����������
+=W<NJI�2=ԙs����y�٧�������D��@��FA����W�E��tO�}����Q֌ho����}���9��?o�a�(�ފŶL`��5e\�٨XP` [c��	s�)�o�Ӳ�ħ��ͮ5�a��=4�-+��B4�N�/�~��/f�~�2\��M$oh'�$uB2�P3��^f�y��15$��0WQ�� ��Cs��
���b\�𺎱�������C�U�	9\�\��T�.���`�����̄��B��0�F�J��
�?�I��+ۮ��u�.x+Yb�pӻb>�(����4��q�f�����4�j�B�Q�L�*�*h���]MPa����J[l%;���=��'���?R�JՈ�U��H�3�x`F3~���e�M"��	<l<
TW�-�'׮�7�����!�&A��PѺ�,kR��"n�j�"�����C)eI�r��!�3��x�Z'ջI��e�2�oW�>�.���2�8Iwn#�&'�i����#�f¥�A��י9Z���� �F�s�}8����]���[��$��Z�&
<���}O��\�9����u쓷ߵa61�F�h�(�F�p�̀y:��X/v�)�������#�}_�u�+��ubj�Xje쟝'-�y��7B@I����J��f�Ku3JJ�*i��w�%.I����?*㢚�y�U�1�0c1�eٍ�� ܁���lu����		zN�G�1p�/8��c4�/�W��`�uz�,C�����C:u'�Mip�WE�6av��FZ��	�� R�=���~�\���4ñ�+�]+;{õ�0��a]T&Ch��o\�|�F �9]��<|�E쉕Vv"�(^�k��X��N���ӷ��%%��ճx\.T�1y�ė����IИG�n:���|R���4g/�.K��U8~
A"s�ģOa�	��v�E�
��iN�y�A���C�������r;��F��u��Gڢ��z�ö�F�;��29���>��lf2���9��cޟk���˒����]@�ý�4CK�xg����O������~P䪶Y�|��̺���V��ED��g}�V�O�ɻ����\��&�拻YV�n˔\����7J��'՚\��Z�}Vh�#�:��d�U,"��ʯ-�Ӳ��n2��{�~���'�I�-���&��A���`|Z���Wo�(M SR��j���� �z!5ҹdI]�3>�{Di���{X�:(vut�\
��淛"P��"Jfz)��B��[��J47����7�����w�#��~������)����v�E@�ެ�K��u9���*�s��0X��]�V�cwTJ�P1�2��u�~�q�n���u0�<bsS�<�H����5F�dC#���ƹ�����-�8.P�b��6��`��w��B��7C��4�e��>��l��T�Sٙ��@��n0f�WUd�V��q\\�Z&�t�Ɯ�Xq9��;�IPMf0�ٯa�����B���u��O=)J0�9�^F@��{�����(�LZT��Y���v@H�̢U��>e։�����橏Y�|y��{��O�\�,�G���ƅ�R�m/A�ڪ&����H���&�	H���h��rGf���"W�:�=�F�r	7j8��� �{ȯC��k�lHuG|�Ʌ��j� �ճ$;�B|+4��#C�,��8��#��.}� �{c�4�>oO�����|r_��9��=�	k���<���μ!��x���Ђ���I��=������Z��	�6�>��{j��8߬�,D"t�U%y���T���˕�#�*k��"�����r4�CY|.�������w�!�o�e8{���Q ��W[�g�OȔ��}��^�ɵp���Z�&�R�4\�ƵT�ty ����ߣO���Зa��^�u|3��Sy�2"8�&��B��C���zW7��!Zv80S�=w��w�"��F�Y�vŵܻ2�d�H�-��Y� �ܦ}�ܯ��v�xͦ�moeh�89���tHut?��!T �J{��6�4�(�US�|~`����Q�K���*B��cퟚD��>�N�8n������&���O�f�吵[����O�>�%��L�gk�
�5=lO1�� �'�dWb^YS۬��8'�"N��b��-Ig��r��eO_�p0K�7+�a��ޤ�6W�ȶ$��w,x
KI���;_t�_��V7��97·ٍc܎\]^����v;������_��5�t�o"�e6�|u�-�Nʜ)5���i�M`��|�a�:��I��1��� ��Q�� 8#�q��o�T�E�<�b��#�DB�ȼ�g�R�U[���o]ԩ}�N>����G�*���Q}wS*2�����p�A��z����l�<1P6B�jtT���S��t�D�G|����=�����J��s�����ŉ�Oq�e�wq��u�z7��������
m	�7Y!R��9�/�F��l���麕�j�{{	�<}^�CH��K��D��FD^ɧ6+./S:�q'�������ݰ�����?�l�r�4�F�@����8A¾�@�!!�Q�Kq}K��d%ﺴ�����¨w
�M���|������Kl�{�
�S���K/��=�3��x0���k�7-�7�&|a�Ӵ�z8�dtc�EF,�S�i�jΒEtʖ֦?������D������z�����}Y���I�n��'� �v>֎�oq����5��kS4���J��)���_V>�d8��r�F���ĭ��`� atC������ :�*��#a\�< r.���k�.\��n�$��c��(9�a[�#nc�I�ɐj8�����J(���4���dYr3�3��X��K�ek�.��zX�0,ƌz�5p��ѽ�^O�#���v���:�@Sx����A#n�	�uk��9.�Ĵ8�,
KV�]����~�4�T1o�U���+�:
ͧKV(T]�}}j��'EE%qym�a>�[�y&	�H������nbze�/WA��d1�RL��I(���5[oD�0���A�
��?�&��aCtGg�:ܐ�L�U5�q�c�YE�$?�!Jӷc�@���ҷ	�R]k�X��"\n%l0,�M�|hsG}�W_�d$���;��ew��,��p�K[�%���@>ʵb�e����<�˖8�  �������`�qϬ�/�d�E/�*�����x4�}��!��w.h��2�иk�̫�wg��!���)B���6�}w
I�;�XV޵ۍ������" S���� ?��_����T5�����n��g�� ��n�9��~tb��Q���r�%�c 
}"�D�2�7����������+4C���FA�\Z�+�U�ס�'%��{@��b��ܿ�k��{�9��Ѣԑߜث旧���\����W�6av���)��Q�!?�]��y�GXM�mSo�����DU[K�)�V���
�b�2�Cm++&�^�$�/k����x���܇z����[��M�<�p���/�BT�Y�l������ݑD+�
G��;����W�p��%� "�f���*��
�0�^���LۖDU���P�?�^j�����̽�h�lYz�����v�os̹�d�4�������4S���-��w@6a��:������kO��%%��
����Z}����8��[hB�w�M�w������>60��_�Ǎ~Q�G� �٬s�'��d�)%
3��ûT�ba����1�D�'�\��M�ZCc豀�]�����m�����[���²���-&W�c�z�S��omJ�;x}�e��lya������L�hV���9����n�[|�6�x�<�P=uK@���n�7�
hO8�qI NU�ꆝ8����=��O��NK����Z͡u}�����NT���� 7e�)wzO�U" 4i�G��:��fW.<�?��z^�����h���3�/yr
Zuq�[z�`[Q���11y��UM���)W&�\1����gvv�B�FΔ��9(�d8�]̖��:;�?�2���֦���V�&@���j�vv�ɧ���24	��0&Q��fG��`�m"��xD�
�;m9#�,�~K\v-�8�����N� ��#b�F�*mڬ4 y-�����O�쉥:�H�P��ޝ�\��������}�Z�~\�T�"g#'Z��0��-�Kz��k�il�������rY��G��P�)�)$\z+(R��_<]��/����ZvmX�
���X�uyy��܅��3l�	H$/%聊*	�&?�Q�뭌�h������X-ɄȘ�c�:X�T$w�Z��� z��y5( � �v�粫#��Q��8��d��3�����]y !���3�B}�E�$�k%C��d,�mU$=+�n�:�_�x�=nzB`+�AW����X'�QW��;�U�eJNf;H�2c��Y�I3����Su
e�Q��_q���\D�9�"+�ALk!������ ů�S�����ڡ��)|U	�5����$��ߘ47������,�\��"�8������F��F$�x;/�(+�_�����i�P��lj5>��`F��GZ]�nW��<94����@^n�H���XҭB�m��0��jS{�1K�}����Xz��[�t��2�6η�c�����W��P���Xuɾ�2i4��6M�%�\�����lc�d�t�e�\(�;���k(��be� �n48K�&�U<K��!3��RK�L�㗙*�\˝�r���u��t�~��쏤I��by�Ngx\>0+�Y�uX:���SxD�Z�rc���kkF���	��M��J�����`�K��Θ�V�>�pL��2^��p:�l�;����!�v0V� �-��� }���:�-�Z|����Z�N����V�h��(j���Sԫ���;�ƴ��u=3���oyh���d�g���8C����.kVM���	K�S�Ȋ��Pj�l���r���]TQ����-m�Q�!$|ƥU�RQ&?��V���!ˇX�w��`S�fHrx�U�o2%��a��װ!ހ�Q��NWj�!L0Ҍ*՚���qխiAr�-ک����hqIphn�a��8��*�D�3�ddMwkn��&��։��|��ծ`�u��O�ߠ�����M%W������+(A-��iD�}���6�^d�&�E(u�Dy}��@}ghQ���:;靋�X����\�,�d8�Id펋�T�΄�� �ͼ*�e��ɇ��P��,�9\��Vp�_B=/�{�U����i��|bK��
�St��G�;�"?_j���(���%���_�
���3i�8 ��ge� �/���Ql���7��r�����C$|l�UA�kߚ���!��G��	�ƙB@pŽˢb���1@�C`"�/hS�q�|R���s��ގI!���dF�c�n;�[ dϭiYN���^��嘤O�V�A��"��:w�:m�ܑi.�����=�Qy �?��kj���Q�DU�������x��x��M/���u���k��K��AZj#��\%_v[S��ivH�������lpitNN�n}X����5���M��s ��b�lQ1W��r�+���x\^����v�Xbk7h־,�e�2�`���Eƙ��q�aϜ��"6-��&iv�ߚ�E��^#�AK��(ko6��Sm`eh_����n�(mW����3$�P�g���hk��������~�!X��j�_`
�7<x�����m�(�~�lc�`���l�Cf:0���`ԡQy�8�"3����m�F�����"C�&ݼ����SId��c�50���6M�g�wR�'4��a����-T^
l�vU-���>5s�D^�4�1�-	a^_���\�*�.|��]���5V$q�X��*Q�pD��:&����jw�J��<�5t�\���gC]�PT:��W�ic�hTWB���@�4?����B)���.b<�vC�珙�wM�w"L�|�Ճ�@�7L�p�䯹�4�A/����������SA;�����XR�����i���Rn�W