-- (C) 2001-2016 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
nv8ljkyWJKiTwdqx4mkRjqccyeMOQ40LnWoF1x5aTpLuX3Zd81PGGrlyEukAsPUv4F7DUXPANOU8
//bvMhib6Eg/LHBm5XUcMZaVPT2Jm8p4cC8hSCKsyBIhW0HNtpxS/qoR4RIrzrVwnNiYhUAJQPQf
fvkWH34MGmkFBGNQd5UETsoxKF65alizy13JxcjG8mNyf8UHGIuZ3jFw9vWMFkNOPeOY2rEW9gGc
TgAnX99oHNyLGvJB+AWKKfcbQ9Pj668RUiX1tAjYedYblqE0xrOxloxmQ815pWRxsK81sRAdIh/E
ir3MNTRe3ZAaGxjjkhpkg64ffCE+iIilrqtxaQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 14704)
`protect data_block
li6P16SFqGhfN+BOgyj5sRR3H+FMlmi7iiJ5HYEkljSsTEG5xq8COjfVka2MLAANO+xsnsWGKAsr
uxGBLFTvoQbz6Ad1l/5GICmfnts3XgsQJv9HgOuojff3802EKLlsupNNJLJPHpEMPOggyR+KyK8J
u1DsKBnNnvGHvZ8ShMBlob0/7WKGEG93xebr8tQJmlH1GfTa6Ghy0WER88lU6yI+WjiimrnXKJ2H
WscIdBjfnDgwW3g6tlZVc8BDqKWiZCFc5wC/CuJlLCeAaQDPj4foZuzFbXsc6fyqHuPTf66iuS+v
ubTy2bUpN0GsPX9SkECeoicwohABTJ9+mRql5hoHxA49Ai0Lcalhr5t+ufuW9XRNVVzP0lwx6qhF
0EK9nBkUBvmxFw5Rr97IzUZUBj6InW7Zhd4lbUsIwCoxTGgVe7qMi4E9LqrHd8PNZjsWEdOXZD1M
FpR8/xUtEDBcYV2o4IlmoDwY3frNrTUUlmmW4lx8AKApT5EB6iFAWE4q7FNviTD2Q4lrjzoB43pf
ZeERMf1bY6Xo84Ydln6lMvUXd0cucgVkneSn7/WsJM7jx816UuRL5tTzKcJljkKxQ63TQCwUgulS
a9uEtEC7lDsHmPQleah+LpoHeECgQtmp1kc82xcnWP5Zkx6CPUzonDqUCRBWOMxfgqT82TPN/9NF
cq6VsgsC6wgWodqWWw0SNBK6sVBhm5GnQSp4e9vDd1W5mDpbHGs5BucQsCABCYiRiFcBHeOfg84l
xlj8VG7voy2reG/99CS6+/xUrjmNv7DA1rLMpQlY+nM8g9yo/8GQB6323bKizQfPCCknpzqXNC9I
GbsfzhVsheU7RsUPfDg9mqC2a2yUfITiBURcuAVg+/WSHnTXOL+DsSl9LmxqGijA6/szpG4kX231
CpLWaYL8kdV+ezaXZUnyVhdmgd0FxMZibkTX4zsgSy7auycaTSbrHWstd3RpuVzkpXR0jqbMd5vU
sXp683P246tRV3AR/+Q2p1NHQr7lJ7AkBLZcGFwYpMA5s3dQN8Y81YcqB1cQYLkTTgUnO69gsIxL
oSWL0EHjUBFT/JNBo3jgNAl9Kj1d+sIiFbog+aF3Avr8EMSYXmnWOo5B1yvya8Wu5tqYB9EWBaPf
T+ksbHrfCRusv4Q+BoCUJOLt4Xxe+7PRMvdvH8daGWXIONARe0acpuwCb8/Dptb03ZIyhavu58xQ
HUXGpFNlyJxuHSRXVP6vEPnOBeCD8opIuEbITl0UsB8CycX9dt4GeCtf+fnTJ8Q8JRqQrafRUprP
Ec/aSLoW3IlJU3+vUANTivEswSkv3cGKKwj2/xQjQl8xNDACE0ywDYpVv5MNM2RbfVC0/H4PgWG9
oJAOW3DbNeEgQlfyigEUfPk0Gs7pvdmshRkZbYERSQ6++dLIzUCepfYivMoy/ggQ/AB1g6w1P/4G
M8Rl8ehJzvdOQXZHtwOW3KfZ6xlQPaW8Qvq7BqQ6JH0kfV6WV06QlWMZtveF2Ve3ug9eJKBWA2+c
WcCTuQFfN64LC9JtTgvHso6nvWg6QOWbqmHvyHhGl7zdRocToI/bemq52j4/Do7H+6T/nvqsgcat
TU0FogoX1GGc7AAm+w+4xlpQY+xsknS1cMPQDGj5IPOvgu5owhd1wt5fwibl6k1qQ93DR1kShcSa
wM4JiKRBmIWgfvbZ7wrnMDly1WkHRAAY7ClQ14uvbLPBIyQ66rCANIYk4skJq8gX1dLJUvvxVUmp
xkvHq8u0TPftyYcvPmLFDhBQhrOVm8v0zpqz7/hexdyjsinD1rfTJKINXkJZziPV3n4FZ/zjZ891
b8NkMzWkztRNJ1tWrdHBWjeesRxE4htMGtEAMidiAMDCgcNLIHQ5JHknJdbZkKcs55bfCMlTBWic
mM/LDR09ZF/hlCB0537hcfuHOGdKgXLb68hCLgORQ0PKH9QxUK69CVGjZhccD+jOg+/OKQ314w7x
0apI+Nd2VDr5oFrOnf5C02JbuMcmdpQVfr5lE43GiPKBuf9skT+bmVPUv5VQZUpEKMyX0eq2iW64
tc6IsO6wORMww0Z92m1/3mi+fjk9XTG1sEwLWuMjnvGGsHWOSXzdQTIR524Z3I+5DVNFDBT4nyAO
Mf8bCSGaORZjXgNIOluxp1iOJq5Z/w3NZ1mBPm/374Fw5l/s63WZYL4PaRorpNYVy95VD3YuV4bK
tIfJ/LSMC5Xz7+UejCjnc3ottkBLqFSKCwHnH6Q5JMGXj2NAhhT+LFIsU+vgdDMqg5XnsmIH+v8R
mtpEzHCMjkSnwNcjc4z6UoQxRUCQiDnIMONwmwZ1LrwnuBD1c5PgaRZ+rfu7fdTE1dLB5tzdzmhY
6BO4Ll+OPxUDNW7Z82M/sDR6hmRqVFnr9twc/FtGP5Mdu9UVbUoAM8D4ooDuM3gklL7UYpyHd/5X
wXzu/E65At48a/lMckc3KWvXDeoiI9Wx0NrAC+vbeKmTis6U7jcQxgwyhA9lNrQrAM7beIUySJiO
6KKbdaK8ldzAk98IswNEzquIRu6H409H0QwxokaOiNlN03CZ+e9dNSUZ6y3MClg31HntLrIe5AMl
PO/tn/r2NcvyQzfXO+2bvHe1UawI9TV/wgu6yDtURRd49hR4ZIPlJtdEJGd+C0/ibrz3gx65rVsc
+j2TJWQoTTDWgZamaW+8ZW3Qn7El/kilmznNeqd2y/sWP3jZON9c0/51eYq6bzwo4EbZUsSdNVCs
IoieUlL+cxfsaD9PJjnmNmxqvZsqwrUFo36QcCmt58atPeqa+RFZ76oNaMM4JPa+nQ599AwD3vFQ
Qx8dA/9jI4q5kFrPsrrnUfZpLvuKJgmHmePDuh2wVSjIO17uamnj5y6FOWAMoeoK/UBSAxJdhn2p
P6X4uOJPehLL9AIedYgv9iLIKdgnS+qhfYyHj8tMZMybCNFdRjTCaKsJSP5iLXKE+AT64wE4fknh
pcuKTL1045Ao9krKLSOiLqMSJNnS21u/q4cTWP4L1QscVLFoQAB9Siobye8EWTbldJh1HDlsoXOd
nP6elvnMR6PyYHtx18TD+Rp4+TUYPz/aGTQ9Im0lTf/m/RnGFcBLhxneS5IkD2C3tnRUVQI9brn5
Utz5pGOY+/ASt084YTSpXogy/VaDgVgk6oLvRNjgapamLHg1immefWKdSYYSrlpQR9L6SoDcvq2q
ra7dHp98FUDdlvOdi3RM/g5jXLnZ7s9Tc4B4/jCry89fmmz/TmXjg/RBlZUlPIlIb3x7nWr4voVd
8BtKQr4CLLuqZuB1IJfBSJgWx2DXGlS3IH5ocM4KTfhILC4dILGynbb7Lo7c5wtwiaswGjeWB8ck
ivNcxFMiwRc/sDT8GOhnf0+EZlmHlPHpaxXk3JWFF99R8i/DMVKTq1Be/c01GlmJ3LQZuqVJqqLQ
HJs+GA/1ScP9IzAdFcIKyXBB4rEhfVfyAJU7WSVyk11gjV7hl2/Ec4w82nh5vy6LsvhkiETLBm7J
t1uOmKgRrQxze5aZbvm2l0INviqmz778TFDuSZ56P93pWe1W1Xn20yVrJAJRw7kX3ZBQAlnL0jDe
X7b++4TFeV0h3You/1P3RAPlzi9/92Sp+qQArexgmDNekjYnGtJyKPRXDkFQUNYXnaS0XxzdDDHt
mSVUy5d47XOO/n/cdcNyONw+Tr7BqTeqAofLcPYJblaoWb7SkX/3aEjyLEkjg4Clo3lZ+wR//xB9
VibfvxQQ0e6Pls9VL+lSCWPx7Y9yGTWLZ5sGiE5aJai9FADv08Btz78kmE+D6+LumOuEH6HhWIsf
v/iKbWNExH4c2DpfJzeYGQlc4OtxI9E5oNMJsZc8e86Zx9m1yydkHP1GjN22Xrz8eHCadw7sCtj0
29bBdVO8c+5XwzsS/sXwa4COkp8DOUyhIhZXOiGmRDQC8vNumdC23SrAIaRashmpTWJYjuug0zVW
6TMYJYmOfcDuZoZsglZliY4ZMi0BKlLzIJ1pKMqPho5fPqMCESwhTTsuFJHArST7jBnuZVbWheQ4
SPfDXnq+7NOiJ5wTrIC7EO4LauzrjKf6LH1zk4xfo2fUZd44nrl+odJGQS+bLCtrw3qQla3+nAKE
UOspqOKXDUVh7lDD9QrI31QtkvGN45BXkz9o0CYU4pBPUGTf3yS+mG5dOS4tEEmwv1sgKvDaHG1G
nanN05nREJ7n++jxcolkABAlAb+lR3SACuS3XFigX4MoB/ZYs79w0xeump4WnIw1nIqmUWTHlxcq
JQlLNpPccsNUHzbuKdTIcIqMGzsTUMNEsn2DwPuNqSXfc05mIrZ7I49JFSELNEUlFDqXM7d1fxVo
lrV14sjlpkYbJOl4mt/ocHhmElaQ7Hua5eItOSIbSbhQ0a9kvq9OBQ8j1mClv0L38wOXTbscx0rJ
yIimGdnp91SR5Q3tiOpJyFQifyl44joNYq2JhgPnZp+BjOz61Ro6jzLYBf9zLdRG1iTAgdkodWZq
36wjH03tH+l9QH5GGjdt7lcDtIjGl+Asfcls60pD1Z1kHKIMMW9g8IoB0Bc149h/0P6NxynlPMaA
vEoQgddR1BIPruYwPSVbgEx4UolSfVtOFwKCi58qNYSJeOTmHS6NeSgvoDVdfEoM4onbTRxH2TEm
MOL9HxJbXr8+KD0o2IqYbPowN7R0juRinqRgfcdKKQHN3AQPixDW7QSnilmt2XZ0n0Lr9KJcAYmC
C4VTwTess+0Habi8QwzIRZFKg7+Ixym6BWTuidk8V867vjHQrsTXutT9SyTLYoKue9xw1dBfvyHA
Y9cW0jitu1oliM0kTO9pyoTn3FmZuH9gfgfJs97quvyfkMLIl6YAjySpI+Mgyt0nmGbeHoKJgXcF
1eemFz+YS2rWswY4mtvZVwtzRdKFG5PUQ9Ha2xQhCFuceg0M2KXBsuIkw2CcuD/3TjvXBaFmfFhV
KLV8XTesJJra13tNzKSSHfV7rmXFMyUAcDzj9rSCa6Pg1zHnfLBitRyId62Mvpy9OgB7pFAz9m8v
ykyaxAFteeFMP0xpxwjiPiKlPMTqAiphbQAyNMIsULuUkfZuaOZlk6mEdhRdH3jeRTeLb8RDyPWx
PpCJs+qimoU09qQo0WaOwRMDqJwPnieGCp+yktVPPlGwrtuA+0ZPUlx+d4gulDO7P75CEcdPsWIf
eBAfgdhGqzMqsAPAEq5lIfTcBABtHdcqMqVtqmbpHTF8EUdAe8p11uIaLGfCiuHbEqa2uMJHRx3j
ZDLa+ArjXOcnTkhaXQvZQr3xJ3+jZ1Y+uc49cGrkKa4+zChhVU8kUXos/8Gb5U/cTO5nFaXgqpDH
qP1jiLkMXjDRDLCn383DPOJye02rTB9zfrYRJBBenQeSMLoUQEJZFF+1cDFcCkHLoKrmgP+etQ+z
xjUmw60XZYFgNMNe4bk0OB3Q3zR4oG6mNaQgtfw/W2U1+kt2ZmNOpTflC49fX4Bkal3iWXgLIn+8
bJ9tLWExPvqlxncALX1uOlINvP+J//klU+rUO25aoaZ8pD5VX6GmXT9IFiH236m4Tuaf6AQgiQpq
5GicfVSPXeGi82AcQ2MfLf6C9zpHFTXPYHgC/aG/Hx701oKStrrP628qjc3S3+5hFr2VKmSwNKvt
fh36Er0w/q5+z3R0g9N8zavHx0b645pJyTnOATQI2KwYx04qZgzHfnDhi/SGgAw0pZ4/NHKFuj7M
Egl8ETvKdK902TgwvO/PyzZ75dQzDFAwm/WNIWi1xOZDPg1APf0g4sdZoQugQHZQMa8V2dmJ1Ror
YV8w7KTuwQdHYW9u0h005B46y3vd2xe1eQygH4CmElwD3HCgaLmCi1ydAZJcPuh4+60fUSspRwV1
rTJqYqQbrk/fd6TDSEfahJBl7/kO7DHPfsaCU3245cgwcqn8Yehe4OCwf5zzTlBEZbNUxAJYJfqB
z1UYb5+Ki9v15KB9DeRTKyvjT7W4CUs2BplSC3ZXFa8uob1O0HxfTVyhdWm4/S9bc6xiPgO+cEsM
WQmuyWOHJb1Fkw5TrTCcQbkXumC6KdfhENWaLR8UZZA79eCdpEgv0aw77/ChRRRq8QLPna6vIoSL
ehAQFDXiunw98zvVqOCLHZK0FXELzru0li9RsdcsxGM6BhIToI5k/m+XbhCm8nlzKJ2dO77daY4s
4qzXHNcl/HuavbUGsoLMvFoMk4kN43okKo189ABM6ILR3IJnlQPe1y0qczvTizUyP9WO9jUfCv1b
ggOglMK/hJZ1mWKOYAJl6Slw4xO6zCsyvWZLmbKZ4oPIOqerKvZHpDx1ABkAtJF26gtItRKaWX1Z
oW0/Xfz5rjqFoq7mL+DvclMswFkyr62hKw5rl8S64b6KmY7bXWtZZwuoNt5QOXsepcWJa5cXH4Cx
nmxVBxsuK6iMNp2RxjNp564PttMZaPnbpdnZJB4+I4m9LLDLA0YnmuXe71590UgeoZKa88ZqGECN
nY4Yu0feyx5rY/ZwKU2e1a8GuDjDQuYUijQQugpvQHI+c2QUbY53bdgGeSK+UJf4qjPvcv5J/EKF
ulUs82tNg1Bq9u7QHaOR4QMQj3HyBWS+x/0P0zsFkLyBy+bGyM7/mOL6GtV9CRIAEAvqp2my9fKH
GbBVjZPmVQSdoUVzqj8BaPNnE7nNrJfbipkuUiMi+1srA/VRELfmYKEPH4XB9eGBMnl+Ml2KvLIa
ac4ROvXjpickFR+m6RpOOnj80KyXdnfjHqKKEKo92eBZICGWvRe59omY7GReMbWhhcn30BOuk/TC
hQ2uZg3KxmpLcXgt6AyPW/F/hLojAzIfFcPExJzxH6CPaWIg5Nx+WMJ3MhrB8d2bdjpNWt6DwFfk
LD8y6f6vnKCpyrr5zfnnroggpr1Cg1rxVrefFi4VWFhmPM8PTB/TNcMhuUb/gZPHVAeddbhPfjzG
8ftIhQCAJOfSthzf+Q4wk0tOGYWXQS0lAdPPSRWv2NzDYm2xDqWqTtv9d8UMHpV/RWO+vhsV+bwS
9ya+/j92rM2OojoVAKPn3PGZwl/bl8oXvEdwcBFqeULnnrfdjZUDqIJPkrHZgUL6YjqEzHDK58/h
eY+2RgUtkDB0rvClMH+A8jw86jvzANnRkqOGxqGV8/3tBYtLBc7MuK/jB97w5FFd67jRUwqgQQxI
MpFB69sCbEw1iFUbPmUZdcJqF0Jy01gDbb6hOQvOTHneDYeZeFjEdW7O0+AhdhR3Ha5wOu6EY6p4
q+DgWPRlmjdOCSpcOvCiLdzd7vpnNChJ9gT1V4AXpBcce44zKKl5i0SBt8zRQu1aUZUrTeGXBRQb
+PFt6L/fgCF0ghFZk2KahNLP5+tOVPHauJ81gm7fd5E+aZQ/YVjAnXIlazLEDD5+7FMshMef4+MY
rKCEOnedQiMdLHvS5f9UOyK7DRd5ZMdAUukoW5U2A8Z0e+cKyXjFeWSRAZFiQY14jvCY4sCIRZ5G
CgnbWO7fF1xBVLMZqWlGiZuBTEV6FBGacqTyzBI4BEUgCXKmf+/+DB0JUjf/x1c/pBdJEbH1HDPd
uPhpYWA/rlsTyJmIedgammlB0mMIA95ta3a6L9bcXX4L/Wm+3ysVrICvTQ1VWOYYaY9ZzdzqX+GX
DEFu2zmmWRK42DKeRVu4wTbXC3hzfW4SMbCoFpVwgE5FsnBeUItOlku+37qQMkkTyjZatIw5tlh/
2t3vBsJGmxroxt/cw3SDL52QKhG+N3UCJz1q4/5bgiPURdpoC+56j0dBMo3qFKrjGnBdLCUygnxC
qsZ2LKCVNMuec/ylqZW2Zaah9dcK2moapQDO9ZezBq99stvPwUglNyUUfu/sgMpUjvNhYL56OWMP
6lEvWkWMwW4UeQyGxJkER113vul0VEb5N8ilhB2/8G+GpRMTBSkwtzwGnPoseNwj3U6X/0zmcw50
hKBYh1LS7fIHgdkDJHBJ/0gPC6AovHgljdp5Shwj+nBVRNO+2Q2CWTCD/WWRjM+ghKb7xJfkp/5n
xJqbMPzEnShOs1pq9/D2PwDBeq7GKDslDXBtgPDAk/2a3Qh65DsM1HUHSBnST2IULwwgmStuZMZy
GIknnS9i4EAzpzY25XYXdmuOX1jDAioSKsX3y0dIAv+1gYrny/LqGovAblb9Vtbnq1Bg8ZyA3VCS
5Zc4YcqhS9WttpG6gLSe9j58odyIJh740fpy/x5c15tPley5m+c8k+metIgS3mDZImezUy2ZfcW8
ukha1TM3x0uKCG/zpUTrgUp3IGNua6xKTZgLFQdzr2OTUb4teESU4zGUMDhR7bmF0bI4YAeX4aZF
kp3cnPaji6mt7lA+w3yw3oOTllXezG03xla2UlMiFk8cP44jr6Yxt+pd6d4fZV7tSh8pRJH0bj93
XcYNjd/62tfhwMYj9jmBvH89RrLGvgo9rI2O6c6muDfegSE2Fzttzuui5HlOYlsuPgm2hP9yxUuU
gMeATg+2bDKFw+gmFmPf+g/iqrFAsnvvhwYV44EI63X9LZDUx2lz4IO6FXP5SmKbzPYuEbqwzQU+
A5Ba3/g9K6ngpGcYQBpTnlCUNM6UCc2uE6rQ8QNxi0v7bMkvYNNgcTIFXOWMOuM49BHxvSMSfhu9
X+4aXT/iwGHSuq79h7Y7rQL9lC7XgMnwybzFqE+lGcODIUQJBkhIcJqPdpQ/dzGxa9mDvtBFyhkR
O30kWWtskt2fPYUmqjefspy4hcg6CI8fIKRUM7vTGOF+H8CdE4LJiMmbN4q/W+Lg5/LBTQKJF8aw
FsiEaJ7XLIvn8CLBhE97odnTfeEER4hPK0BfsEhZCy0EjnEwHphhd2GKEEPVXgPfiobWq4Lo+oZO
C3+Lw7xEhJ1NM1nnx9GOqIHFTPrt52m4CE6IsLgCoGXudHP8b1OOqJTF724CHvG3ohtkEJKp7m/6
N/TjiRatEOp4pSPbL+2XLSBIM0+FAvB/ze/qTjB9OYbvrQw+8gH/Uo/xCW+KHt1TDkAm1wUUR2fV
avlQEZcSkc9WBJwWSEkbjkD3rtjX2S3gFQIsBMqBNgxcPTE91uXAe1BrC3waGgaJDCej0HfBs3zN
+XU9afTFMbuPaOYdjYUjHoGRBP21+n6o6a5KTXqYKfiIheYTWdxL/JuxwdbgrZUjzTf2YAZr8Wk0
PWlR2+Gyv5wwvjOagqK3uPFBp0ua9NIgqyLyAwaNoP53xKaGA/M5ONWKt/Ic/k525RwmQJYHkur+
1NxhReyO83OdPooI+0jz+Gyl86rqmVJDG0ZH3Zjt2F4P40Tv2gUJsiC1zIejiBfpGV1m2gyA/i0f
wg6+z0ujG0Mgd1WIWwE8L/XXCRGEk86eUxTsGBw7jgLMzesyDTAX997XNhEm5iWqaF3XviWkjPr6
o+hLW9WpmF09bWxHSmZSnIn3reJJcJEepdKcqNl5cMNikIDDAv/mYfIOMu2NpYHuCBbIsepMbe5+
PXhAWRO+lewS3Bn8XQFlPPmMVsnSr7/SY4kLrBTLN7s/EUljNHXnViSg3e1+ZpkmOqQUbG1YSK75
ioiv98nwFBryF3FkBUNFqT66/SIQzSybUBHeA7GBKp3hjyZEiMVgxX7DI8xg2InnUfsnkO0QDy9i
PhP3DAmDB6suKjMV/eb9WwJeKot2/lTS0nQ+ooCpLrkWmwMYrntwJln/JXT2qrAfQ2K5Ggxl3Lqg
KEGi9bV0IH9NKqPTKn/YpKhHrKDZf+V6Cq3cghaT2yaj9+MxccZEIhGouwH3LtfxfbJ0pNAnv5DK
gzTGGI/fChJJZajJlvNLHQN7DsjibFlRZ5anuhf8ry17lohwJzyi3PNivRlkojql2J/vZb7J457a
nr4IX929yiJCbjg7AwmpxvdDnL6oEtcgwl3T0BcWMwS3XWrw6+pfS1Vor2T/4YUeOdoaEDTUSERl
0qzveE5U7R/DjJqnsLExpicWQ+525crkx1nrGUa0H+ogT1M9mLeu4pzhQRfycHQAGtmaP0cNBuZS
j+D81AHJ4kaBTEtSeLuRrIX5yBZXDEDtKzjG6VjdPh90T2qTs4vwGZWPWyLkik5FJ61BRnFgoQWC
VNB9Loko6scljVRbUGDB3Mf+Nvpb9oc9bySznvMqqFIFR9tX4+Kv/n87RmGNgOsQnI0Ulmft7eYO
P828mgp6QpNjYeYm4WCbQiV4yCSZN3Pkfqeia4QPLsiJpT3Cye9lWMyYDyAfDySUEqotAIbBSAe/
+aSCYLlOXno0Z1vipdiKQIs0V5viDWmht0gGx8aGv6SYCdVgV+VxugbxjsPj7Zt0/qOnfURbr+XU
SDZkJpqc77+OCPdC3qUifjCOiCfXEqB2QQzdoA0fFSceYNASGn4bRrx2rMmXbkvSEGDs1xpOuTDx
zNbVc9IgcazPKRUfe/6iElXS4L5cUFEEruoeL0ejGaqVdjqvQH/Dgt4VFu8FG1h9MOhiYi1fQLdb
EnjTXU4vw1KNmdZty5aBpETk6IXDpA1uRvtmfkMzem2+ca2J05gWe/t0GBXIcgLqMaOiU4O+5d57
4fcQLt5Zr8tOx03z5DKDPurAFXjt0f1WhYqe1Y3iv/ZMnx2qH3tAjD7nlfe4AZaSBA3Bggzz+NaU
RehB9ERDZT5sM/HxvTsOHBZ4bCEPULOP+03uunCJfmszCbJvrvTPVxvCN4I71GVRkg21oScssZBx
k23IfR57WMuwYDMNyVg0cPvMlYumt8zHQrQhN0qDAjaLzqmBe8UvBBvsRxV2sbktwOwh2tJJA2eA
n0tDu6Bi4eHieXwaeZYo/A0cUeNOi7KUeoczpfV5JBtseqMi/nMcU0cCjDomhyUuasPOuBLl5gYy
qk7O4iJDZrZsxKrHxgoCXEhUF9RmIUFmn2YrVgcifhYeILMOogUQvKHhIKSqE1BcLudMR8eLDz2E
fObCMnzzLNjfkIYMcjTs5AMnCiK1ATJcnDm+zyeDD7k5YMq3QfZjUUDvfMTSjyOGuTb3y9hVbR8k
0oB/kpq7pPxdw3ealBXgm3MCf4053hlTo7WDyLiHFU7Y336oiRSgvrYixJac1VVQ+YHu4bdXBH2w
tu/xWGdSkGeFO3jgdRf2q8pyvPJPUAozvoyJ98ea5vWeV9kZ7u8RieegVmyOSHR2bOyw+3vPEjL3
QMzlzkr9LZgYmXKXn7AZVr7bCDNKS5LgB0uf237msj4cPlrTs6KeTsS43nK0+5Xb7SN3QRc+FmcD
AN3e7dKWttcYBMVw7Z/9MpLnT2gT6uTbuJ6SMDqlMwXN3EPDXfw9iVTZWFNzUpvgqdm7atysOsa8
gG4UBrqHbryQrWo5xfIF6D6B1UM3Ouh0Efx+bbCav4iGzAbzlaGTVG1d54fGn0SnEoFcCAWYwqbq
ABKXbStb9Ak+UC1x41ktx5e8yqal3DFQPjGC59fKd4IiaK/7TIcYikJTlbT73hGTFfLqS/BxHuTF
hpW5uO/771PtnDpL8AH6ZN2ol3TMwA173ZLrAOq+9jF+GaF30SjsH48DJ1U3HlrxA/ANpF77dmbv
GN7qexYSKCwkWFxsSJsQteHjvb+tZhJKv1vhVEIyfCI6ny91W63G2XrLlS1nJpo6vuLskeC/fCK/
C6eLGymx09/56ACXwwRgEidVL8cWO5eCrQ1O6PtB0Av6aaezJXew8XzgqisiYyclkRzUKLnZ2pbE
C95vvPvstuQTgbgzT4gkWJYZkphDFZiwKvy+GUCB/g40aseCWca+6dsYtqpvhYry44gKEOntLOCe
6jg+osG/0hU12v3m0dy0fXy/51H/OnL12qiY6GRbWzJwgt3NVlnGF2ZeCXQ67YA0EGDPqguSLn/O
Ooxs/vSWBaDuP73Xzc6Dhxya+qnE6s6EIkUBFW5/vmpTKVadYY0NvMXqJXNodJZYCO9+A9d5r/0P
dpyVfkVUzCtFB8gBcdJdHHTu2AnWF+bUs9UQZYCb+3i61n1x/VjUpfE8k7o95uyuDUC7AehKaRIW
JzW6U+AzxtHY6IzQ6byRI7LVL1fyXRT4Ui5zCkMe5EXHsoGSjivEhLeQRmN/cPwp0s3ubMHv1URb
r6yeNzkNQcwk9K8uFdW1KP13UwBoSAWztWrr6S4KWqG+32hyQChLylx6RscQgTnBPHsG4bHA3YHP
L3MeDEFXEEHQfx7so/d+3ITJRl87nRgKbfhxWl9ZWpWID+Z979VBd+kLP8qHWMnS0daIL/kzVKKY
MvplvIO0DE8TLmOBHqyKCJmpEz0KKSwYzUD+pE8KUIZ5873BVZynreLZ0YJJPTeVbhaFKD4PanKi
CqfH6f+HFMg/7ZVNurq7e7UZcaK7MVYUB0yaUXDlL3apN2hcSeusgbUsPNm7P/ocFgv0xPj4e5GE
YS3GNElNe9pAzF+lYgUOLi1EzfmCE1XVZV6tTpCvUD/l6RMcpZZxWce6gVWYgUTmVp+brfAW36oP
tHaIFy7RaVAfZj59fF7zUVMhlCq8QZ4/c9JK4hROOaelBwu8t6/YIj3uxPOaLEksjqDQobuKsDiw
yNjyfi2vJjEhOfXnVXUCJoIaojFUGi/8H/UGGHVHqECTUKjIXOy5k800MTl2wNcvGM+rWfDXg5Co
pLDSNOhZCYfY9eNzLWfPlFCndjQjYy0Pih2Ioz8dyUDac7lZCrTMdlAgu8hntzBc3fEsRvZbpVLj
y3VtTNJwFAkH4L3sxvlvMX5aIpHDWR7b6uzxDz+4u6SW+YYPojfk0IsUf1/gBTAHcUQ6n8pgKR8S
JSP2MKe4HpmWvrVrxyZZwXPlHx6E9UB0dlMs7HI7E4tp8GioalUipDlHgXtzSVBJNcRpMzbJBjmS
3Q3mJKG8tcrS4g8nFhpzDxc16FGKpe4d5xF540bdCKg82KN3kwOlyHD2PEkYjvxZFGtP1JPfQyfX
iznsISFgDwdz35HW/iPuVYlvhbUimdpAGWJwl7jxsIZMO7gpcOENwJEx8ll5n0j6/3yTBP73I4Ke
wzvFGkFSYrrdHQv5Ey09iE3cu3US4iBMyEA8iMgsYBA/09Mu59SL2B22KkbVnNlRM4+xDSxpsYdk
lIQZpvj9+wn2Aw6L3KUdxp1yjpfv0li1kiadXvbpmLOxLbRQY9t8WewKt1cGXOOg3UTzkWPQI0k0
fVo8CXSFzR24wlb/3TnMDETjH8A9TVUuVFKExnFWjGUIyLo8yakAscYD3k6LMNKAAZsDisQc3C3I
jmfT3wiim1z/laRVNnaQIyWGkePdjCcOXmCJcf0hJSE88fqQj37xJqDixBmQ6COcb7MpzO1PFD7P
YUDo1GakXHaossqwagcZQ54O+4/jYg8BOPwznOmBvZEMbmZ9DSvNfKuq5huqg4Ax0xJMxEZ8ey53
jNWnLcQNb5c98jArGu6soJfSQpiYS45bSyC0nwT5Olzxys2TyRW9kybmhvh5Cdueh/LEwbGxAuTT
04jMM/7IZIayiboUIhErLuxF2cn64Q6RDxUBqbt6PR0Uf+yQQhAcSVioNW7OWnFGrqWZTAXlgtyg
jbsrPCBpNWhB0vXgB6tp7EkvSBr8PlvGTpQnLHMFhYbmR7E1jR3O6T+udocypbJfOvNALB7eN1If
pa79sCSHPL+lrdGSiu9060VFNaS5KjaVoLThzDRrEKRh54aiSEMn0HWGkrWi/at44btvgXYL1MoY
oqpMpUbfNADAB7xDRLkEOO6o94BilZbKpOevDxxVaMDYY+8q+X+0KVN0YdVxPXj/B1+EK+nAlI0Y
wa67RivBoFclFhpxKBdXRnNSgc+7qMVFGc6oMSDmKqMxCgVLfXOS2/Kgu3n3AcQoU5sFMSFnwqEb
Q+G0Zi+DdUEgcSddt04dHw8ukVaMu8p4AAy+XYpyrDVGNtWVkIoncNAcwFj0EZR/QiN/1XrPTZOM
UgiZD7Ap5OFj7vtWr+QqaXY1jA3JZgjU2PK4RP4duemtazdfyqZyMNpKrcjhlzefkvei05Vo3nR6
ITEJwP2y58Q6ox7HcSz74PBGNLPsYSLBTkm3Nq1c83tmBTltAiHumjkw8JvZo7MSZobBNwIKVamG
qsslvcW7cUPJPduRj+X/qaPvJDk07TNL9OO3O68/shvZs5rT2Kx8vze4LNVM7ia5NYbPtkgbyGlm
BPYlBXNePyi3VaAvZZXUbjJjHeDN83pVRSdkHYFbWplGAmivSEuJ4fjEDpQ5WMPtmMlP/x8hpvVw
b86VOdtWjpVHlDobmv5hfKkGpJxAj4UhNZ6DI1VzaNO9ORSFBqwpuMIp5iJwnh4ZPYjdqXfwPjfp
76q7usONqJhSBC4mJb5eAGAn2J5x+NgRa+NhwhvGBqIgMsgN7CA+r/ILZm5BW4omC4JJu02VRCN2
eX8YLQPKWV/YmGNDbbuNBB+MUVxqJ8Vz9Dq+fHFdShBMU1rJXlHrZeQys3jW+guKRPGRtL0F4BU6
RdPxsYHLqzIVPiTK9MQof/9lxy8zU3fyKn/J68KzK1oWXtiuT426YUHWA0C/TTef/GPO+liTM/ZS
ppVLENhhX3oP+VMIOi1wGlyMYqtg2U4qCap15vPcvdW67Ng90oxTpLM7OeuqIx+7rFJ0Y1nElOua
1fZly3TOYLn6W4G9pP6dOFWaoFG2DhB/Vr8FYVecngv7J/8tXQEDAI3KUAM6OljepWzTKoQsKPsY
ygWCKIpEXDTaCZoohshDDffpYf8ApRfA+CK5zxNxT0orRaBlJSS+3A/PeWiMkF+vFpWcKSL+IGSz
5FiNz2n20RFfAaHayYJT7vRsehG0qTy2lp1RGF8wbOR3RPzZ4yRJbkQCZei+FxxAXRQoPa9JtZNk
vJISGPQIXs6ReNdTvggsW23/xbPqUHE7okP++lQaAf0tS0ieC9uvDwTqHcnSZv7wmyKRnzHGF1Zz
UxZ77S/T1ZI+6jSthuCnwCoKg8XnC+0oQy7ANufa6DRYSOTelZarSnkMtfaIkJYrgIFnhKFgKskT
3EBHBwS5Vt5N1lXWCBM2FQ80c0CgTBOkX8w0XB1ysQJx9EZV8fM2DsYDV5pAITOdl/cSRK2Tm/SO
c5i5IvqU2SSYUCFfdfglnQcr5XqcHmWrl8Ir/+Z3eiF3zqFg4MiuAuqBB/qPcL0xE3ZxjO2w0B0j
QaCNZoiSkkwONYLvTJyp2DE3kypkk646rPt3bSMYkHIkJxvrcOKFk+Dyhe6f0Eo7Ub3f2Bvoyy6d
6nqkjqbAGjOAu7pkbeeplPaFGt4PjfucC41tT14HQSpnihfyBaPJ9XE/TYbnvXzLvBze8mnSRijW
KVRC9l2TRub1b2EJOh16I3ti6EGuJ/8j8RLVhw5cAzenn0p6ulxohATTrcYTXuMlMZ8/OB/7WXR7
IQbLJirImL3V3uW9JFXx3Gp5nUhjo6Zi17Osxx+fbsoduza3oYXyydQ6ffjjSUOPzfaURgGPHTV/
RC2QplfZHrEQVkxG7hXdPh05lNediYjMPw+1mnSBvuDX5RkBLbB3oy4i2MzIASrkXW9PRJWO2NXP
rkq05IRVHl2BZJHbv7NDMDU1G9tpTi6yId5i/e21dbZAMBFUc398WtiBtoArSFYmECpA/PUiErjD
jJAu/oPK5pcDo1lJoqAvgoMit5eSY5TDzg3M+9Ls2b1UwHCXdTkTF/OCmeCzEoW5ZxHtyGTqGdty
KXMo01++fsBh9Ut9M05jM2bXHhgjiUH1ETqrW3n5jyzjcaAD7efwvZMlRb00XW9F26AAHJuZ1P/0
EmMAg+ERCrcRcguh9rbaPM3SyMr6fEbrz6LTDUaKE45QyTRhsoEkRWyIXVJr6z4vy7Mjg4FetXux
8/C5ppZUHROm87AEJ2X8Cr/WU/v/u6EiiZY6g+UYeLhgCixgzfAAet+WFVFeF0QwfeYmTsdgTn67
Dq6KDulDKC3/QFC5LmLuM1NiigCnbYDjnmDIJQNRrGBfZ2pyOxmyKJXfoTVeDzuVscef6ej1V/ho
3zXXMjaf7zBkCt9AVGH8lVF8Wj2vJANoa86PcFIqMsWjrwqBNRMQp1nG58s3QH5fkeM/szs2g18Z
FUuZXaenCnA4nORLUOYrSPhpJ99H99t+AvoWK3BlWPdlxdy5MhGoB76X8UFcG4erLCp+/mxSi0yE
Bxx5zSnZ5ZYWrahyUUWdj3Uu6X1TgWcfVUNCjnsDEK859QVgokC2E9+vRuFXJQUE27hH3E5wN8wg
WKYG5dsku5zCauIHViBKB9wRUI1c5kAkfAygjmpnL/5xnWEQkypuTzctqdDx7vJg567pJNwRe7qO
0aodUr4ztkO09Tj/xexL4CjJQkwWwj8gV6yEIzm6G2snIOo5SV+OYW1XUf7F7jkKCrLGWt5wcZoU
JUouFObqXo5UCSDFopf5LO0DtS3xtXL9IsbVcYiTkLyqQH+xsziGAm0ltV/fNHYVn7fg+wq97grL
lQA9y6iTnrlqd8trgSnTMVABJIfIoQCYZvUOV8gOJL3ZiMG4GQxjWIHeZdOncVmO7JiBBlrpuTW8
4lU4hOqFSTCzrtxpaGfChV4Apkt3qcz7L7mc7CH7qfDk/6cLwvnEfu9pZ6KsNpUPPRetHMEDnWb1
0uk7H+blrhrtfjfnbUsd0UetuUtKpLXCTg991cx/8NDcPPG/MSofJT2q7ppUage0pxPzUO8AxPPE
etPkSl6xNc8HeNQ6z/BL7xQ3wHECjr2eDHaYuPEWHMMbrof3wdILC43kCyCkPfoDhMfSOsC+xFC1
xEsu2KM7jfgAX7sebdAXIqIgHsMXS8pUQKoZIH7+U3UJJUN47MKAKkjyzxGkssSA8OfeCwuKMRZB
6rT5Gl+Fb+8cyJElSDwrvXn0llRiKuGz9/9NO+Zk6aDTpgKbjynRwivwu1hoEfqq+rn5nXdpLMFw
h/f0BMv7e+f8hl5+2pSQloezKTaWzf9comCkq2Fhf9+8icH0vHeF8A6vwnGcHbVeNXoRiKpK88wS
VlGgxmbc9m8vW62beblCjx1P5opv1Y8mNYu3lPYvAInrfXQy0vYqWZybBIzT286Wq5JkEWD5lluF
BguK7vbKcE9JC4QbE9fQV/RNJ3/wJU9j9kO/3mzV0ZKUDFn4TNGqaYG7EwALP/JN5TlCMB0ttZyR
vk0jNRBA+WBsDAObyylqbsHZnl+D9Vlcpc3OdgdrTl70Ahtbry0NH51bpGYh9v/Acj/ba4/Iyt+1
VSC/+0aKhenLiue6DYQQ4Ix/TuP/HjSSpZosSwN5XWm4LlRjwoAxzUddb556A+jtQA4QB4596ISN
7fOKpMYtqV9IJ967iJ6rO+8lF55N9PWrdxm85lnZ9EM7l0ehb5RglSvkV2cG1jW+3EsiFtJWanKT
31Hgtp7aWCNoIk6n+KHAx0rLTqHa7nJFsSwO4DblUxbx6Eq1fieIU7snd08Mx9YLWV48aNSCuwpZ
Czx31MtcBSFI4g6JMkO4aptyvqS7d/Yivy6DGYVurtFqaf4F34xPDSxlko386434K1lWX7SP6r3U
odlSAL+XbjAKbh4KZbcNP48TnUUiM1QDjlms8e+GMThosCvq3pqSTkwYcOsemfmAPVDRFrmJikiF
gb4K2RjReXcYTYN0q5OzUOqvSX235gHQbroAEymlpkfGtebjtHgq7iOAQPuJXx4kpnsv6ofvNhTA
swXY+oUEyaljM1ff+RzReySvDDNRoYVmapOaTk9vxmgtmznyTBD1eaZ9Fvaqvww1ELWzxoSs+t0r
DBJPvdMWfdP+8jBHJDgcPPHZwMCRNbI6j1b0n+6XboG4TKrTOOVGhI/ujw6W/l77LBP0qJxDoeCE
BXeDimfGezBTOA7AAqkTWPlsy7becLPbC7ip/zUG4K7toYneUk9rXpchb7G0xYquKn1l/uO5jqam
mpR/GVGhB+YY+nmd/TaZHYqPmC/VvRF7rsIpxRa3i5K8vS9BY0w1IdpdIyeoRSGNIpFm7/3373kz
CXsVwrIL0LzYYgKcD+CvQGxQGkhGLDbto3dvpePbh+e2vS0gG+IIXWIrCQM4sB0IYNZit2dWeqM/
rCuHDPsCAC9C4Aq/HAGessWXXUtn/FEvO+ws8izYUPYy2sXtQ4Y7Ninqf4eMyaC9TxMeGX0DjhE+
orI9q8J3UlwEJykWj6QCG9lqxajzakUf/tXw4yMVjv1pL4a4P3fxoEL+2gJ89Y7UoNgz8elhIsLZ
SnjEUcnel2uOaxQvQjP5j9jGG5t/TrBX8qszT1shnhFO6h4y+Gto/UgYyYM495pJXb1PaBVA9RNY
Sm30f346E+k06Ovz87f53EbTYFDZzD/OiYpeLaL2dOVY8yWuiuNqII+0HNHoA1+gKWRXx1oxLwS/
+ph/ROcS/cWiShUSvurUTMIRKgbGJdGGyOROak9fycVwP8imyF9zJo0rEwkyoo4SzcjLyOA50Nji
xf6oGBZDpb0QLOiwOQKmdUeMzVVX6NSUPdbidi6WtN/xYKcB1QtqM2T1zaT/eGTqOzVaTkM+Cgik
SlRwnuRYstoc7gDukpmmSzE2xYMGOnwwbwMlkJ51d7b6ikLcP3XTrHD1wNRH0tWG3boHndnNC4y5
zcVDtiJZyixKC/OWagVpigzg92c1EkXgxSQXXXRqi46bfmV/jx/cSZz7iRksrdgTd/kerBMFLzQP
Pq6nlUFT5gFS7N8bmVr0Y4CLLhm9mm2m/yzEccYkfVOB9EJNZ/OQLCKpxwNJOOue3bPULCuyVISl
Y/RLgS87b5gKzZdr6CFb6UyLL2PTfEfSNSZp+nqdXgV9XV9ZS4qARC5eJrwnmoKIlBBMVTif2zeB
hsafcnUdWFmGIvjNCDz9e6C9TQjisDH5si5l8oS0j8R0uv5x+rxWTTk4chv+fyhR53D2fh8LurML
biDS2O6DANIEI99Ve434zRf+Y+1Ecd3EUGcN3tkEJfZJXIdxT9zzRUJ5PmwBEkSZCvplfKo6vnTY
rCIvJIZoeFBT96cikVI9atQ1Ax8zW61fCUdKb3MVUvfnseFsBnIRa3kmJ5pxln++IJfhEM++otym
kF9WynqmBGA/yPG1keS5rFWTxOAahVs928NGisiArcoQnq3tmxUwOiUHErwihg3aw2uCILgoedAl
2xDX7EwpH2aU1Uxbm7jwbC+koAyJiKb4gJeQnjOMsa2pIsTcwU/k8fL+39nD5jWwtXSXC+FP/bYu
aS14W2AB5HIyBfOqYP9LOGR0cCac3WmXgz8f5Lo6U7mgFRL/fbebB9RwwJW3deTe93dI+elroFD5
8MCXfYzXFybYRC12ObvfLId0vAcMW+Vo4I4GvS6v+Bt5mwwVKL08m/lEOI7RTcsVZmFeNaXlABsN
IP+rXscvlxlpStK9Nklj1oILWowGFSyoqXRSA8l/ikdgDleENL566vBLIMpYUvKS5bOhKtTqIOD1
lnHC/gKS5J47j0yyYHiIWyDA2p/l9/s8p1Hj9YUjnjtJGaIRwyFwv47ZLtzTaOjDF/3xf5KvIwCu
BmZAzgmKsAxBn0MQI7NZtQSqEhLvX8koBRmoWYwdllbqZq0hco2BjwMmdtQpQvXihKqboiJHMqrG
C3SD1DDas3wvR7Vw9eqptGpOWsmUGgnTErz/7pRQ1qJRwNz08eN+baz+Xh7E8b6m5iB12cCrrlwp
PF1XftKhaTv0El3zB91UHOAv+VNXbHU+oYy8h07FwWCi2WoU5fuk7+3Hc3x2ChGTPRu5QV2HIQ==
`protect end_protected
