��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����N~@#�k�0!����+��=L���0�ԴZ�2�Mc���ZO�����=�����վ�	"cqw��a��TS[��{=:�����K��-�մ�(��k��N�-� 偙O��QZ��~rL'�x[�i,mׇp���O�I43��4d�,�H�����SN��d���3���r��m���̨T�I;uj2Y� Er�*p�Q$Gm���p�V�`�2^���,hz�<p��l�Bxt�5��s��\yq���#�@W���f:m��T�	,*�񞭋����_��㧋l�	�\�:��uGd��PǷ��N�I��_����Tuv� ���us�(H�~�{2H�:Zor�Q	#%�3ˠ!��iS��95�,?�.���/�F�i{#���Tp5����Ҥ0{%���2vpn���X�����@l����3dc�ק�3	�Ed&3�ZN O���z��s�yxӡt��v*}ԫy nj#��lc��m戭k[��5)�A#�����8�!�]�Z�s�M���t��w�!��'ÒE�rv��Ϝ�c@<U��\tq+��&|�&X1)C�����r�A~��B�&�����s�:n{p��͠R�X⺂L^��R����c���f��J^?��ܣR�O 1�rV���:��T�4���AD����˩�F�w��)Dm�O�b,�a���1$��c��7t[i2>�ޔ0,S���󧇳Ϟ�ᒨ�-��}�!6��Jyv�醊�^_�(�H�(y^����o#����X��3-�k\8�M�T�"`R�DF6ȕ� �,5�;Ҭ C�k���1\������k�t־9�}���� ���QHF��"��t�9 ?��{E_�7��!����](�S��0�q��w�9��=�i]�1�GʦȪc�W�XC�|�$��}q�6����zf(����լml�dz������*�eLD�*�,�m�]ہ6����D�Gw� �g��' A��)�m���b�����L~�B�3A�/15�s�dm�\��rbY�6�g��x��E����Uf��)
^fd���YaŌF�<���^1!�C;4�i�@��e��f��1GY|\0z��Wea��".��������Q��F}zm̋�{�h OSK�&y�À� Q������e��5.��ѬQ��G�P@��S@fx�f��{���A�������U�ǚb]wT�sS��֬���/�B�'����	bk�U��p����"�-m�U.+X��p������J'I�^�6��?MwZ��ݭ��E=Eu'o�#\t�>A��:Xۋ�G�ӎ�B��7�y�4�)���D���[�$zOy`��E�:�Tc�Ʌ3�.<�݈?ᚢY��n�V1���k��3l� 0�!������`z[�0�P�z-C-	S1����G�F�Q��⊢֣F�
C��\F�]
��/��fb�&"Ƹ;���!�dcr6[��iG<P���b�mmRU�A��vB�ą������#s��J�?Ǖ�^���H�i�b��q�7���� lR4��)���EO�ɪMf�L����bb}D6q��H.�YU��%��[�D�� 
���)�Jy���5�N;4�/?]�q���`��!��2V�b OP����Do�%��YUN�ݱ1Թ�`b���^m�O��-���Z)GM�N�.�viy�� oC0���uQ�#L�3�Ifk-	��Y^xxPx�4:�C�A�"[Vi$���|Kp�������������^�_�S�b��,�I���X�@���ڼZ��y]��g�R��9�y��p���<�7S���&�M��"ti1�Y�_F?ה�-9�t:r+��!G���4#������Լ)��c�04�ã��A�T:�5
����媿�bJx	�A�,���K)�a���ʑ+|�XNmm���$}1����=uD>e��t��O�Ѐd#����9[j�Wjr:6�wNx�����؍:-P��Y��ޢ�y�'�D9��T�
�Q�'���?��zە�h=6T�ga,~EK��h�c���ҏj��oH�S�q�����S�L�\۽Rt�LW�4|�!�*����ko��r>��*u2@�`����{|�˖<���L����h[�q�T#�ai��١B�ս}�j�fT\�\��N�AD�{�����B�����ߊA�{T%Q����i�ؙr��|�1OoL?yp���!pz�J���@0�}�<^�[�
��hQ���e�����:C�̡�p����d8�u�D*���:L4�H��A��v=�:eđ�����譳t
�:�#Y0@�pJ���Ǔ���!�T��0��	"�|R�E�����x�Q\������!��y����5�Yf�m�9�^��z�H�f���t�{�U�����Oֳ�D�����K7��Tp_0'���F��+���E֦~p��uJ��hqw��鐀�^��'6�`�Si���m�vpXAŕ��wR�@˫"��l�K��z�(����u6��Ҡ_Ee����;q�g;�OG� W���A�;��
B�������}V��f}aF�NS�,.cY�p��A�r�G��������=J�ʞ���t�?�B~k)��8�N�C�LR@!J�fz��������pTQl����dK��S�KdF�~��h�O���؍q�p�-��������0�Xh}�{�	�W8��ѪB�@��-���U�q �l�����i.���3�lI������C��ۤ���U�.��xӢT��.��5�u���M�U������r"�����>�+&^8�VH�����޻����wǶ�>��\��q��B�� �����W�iTm|������0���cF,�Y���Eڒ��g֠�K�!p�7u,W�sG�ʘ���1��P�QV����^A�ҋ�d���Ή�j\]VS��8��@݃��1�=)P�r.�88��^�]8�x���?R�9�ck(�]�I�����Bʪ�A�KY��>����24	�o6/�j*������C����G-RK����Bp�U7�j��[Y��p��1!�c}����r�M?A��=KF$�N/�dMJ�?o/_AB�
����3R|{pWA*��Ej9�(��=��k��ɩγW�N�x*���ɰ�=^�p�(��ҍh�%V	>Z�r� ER	�=�ޜ2��Ҽ֞:��Ԋ��Ro�hC�6�+�;q�����:S�����8��f��n������yh Y���p.rf@�f�c�L���̱l��}����E?z�m����g�͸@5�H���'φ�"� �+3"��L�*L�s�SS%t�0?��K�THB�����;��g�i�D	�ņ��*�_��C�e���]"k#)_o��h +		��c�#�Kb 3��gҕ�`q���f�IxOs�J!��ul�U�ʳr��k��?�"��e��r	�������LDv׮�_xәMF�B���ܕ���Ϟ#�$���@����%6���6-_#�|����3ؾ�u"�l;��ǲ�# fS���^�x�0;��i���)�K����Ud͆�S���M�&��i�������V%FJ�������)���G�OZtrk}Q9�$j�<7Ч�^w�֢hF���e�f�YR3���寗�A��Ҧ1	��(s�^Hy�����u/�}��)+�a���q����cSQ4���YV�w�-��w�'q��y�!J�4ҏ[e�6�D�T��@��^�?��1$>Cl���[3ѩ��q«�{*<$��D[���.�毿ZU��n��gYuKD;�R��uO�G2�6?�M�����o��6m�ґ2�&0�KH�+-���N��Mm��F��g��x��?�R�/w�4,"\�>��^v�-,���k�w�Tv�p|�A�E��$�"5ˠ��%���wɦ#�-����p�}�s�MX�& RC��A|a��� �`b�7W7�o�;�u�Q����`	]�N��̝��#-����ݻ[ib0�6����VN:Di������<mZ�d�C��5¼�nc�y}���e��K�\�^%�>��u��w��vɕw���`�h�*�j�#������!Rm��q�_�n\?�a2���zu��a�����ղ��g8yd&���Q���Q�� n���m��j2��������|�����CH&�>�������ˣ�ĩ]oo�RC�chqg���~k��6����V�����<p�9K���wc�����Dh�*"���]W~kt�ƐQj����䏙yz���@p�����=�&�塠
	����=�;:�'�y�zC� =�0,� ȋ�4�2�Ȩ����fJef�+5ӂ�W��N���ߧ�e,��Dӣ�FR��V^��:a���+���lc�����bob<���f2�n��w���j������>Õ��oF�ϼ/s���o���2�ɸ�����FS_��QC�^Ep`6���9���{x_�D�~���C���r�R�P<�����N.��W-�O�Ѡ0��v��x�5ෑ�_^���8x]�Y?-�q�.����Wg���R����rFluY2�}�z���f���R:����e������,҆�ƍ�;����zT�%����|M\�c��,���.~,5��gȏ�GP�&lWE
)�`�$-�@���TS���RQr����O�����d��P�w,.�pgۈAL��)+�V�r~�v#j�fZ�կ�E����������S�����D��#,$�u����i�������;P|5�� ě�AT{��������H��BLt'�х�>ԃ�RJ��XE��v^�0�	h��`K�nVW>?���|�5��hO�@�R<hG���77S�Vf�f�P��˒=4�٧��3)`C3�a.]��K�nN[���c��%r	t�"�&>��`�K�����ü��@,�RS'����a��e�9���>^��Fov�o4��Ŝ*"�PQ�72g �S+�#�H��V�hb�:����_1��E��NH2?"3�=w���ucb`+�L!���LXg��*�T���ĥh�LY�-��%�V������|G�扴@n�lXR��hce����+=���tҏ�}�	7�h��'Q�5����#�C��dVzs;�>�TX���?�~ @�4v{p<�P`X����.JZh� ��{�����Oem�(z�s-��2^���>֜xU �|���E�����R3T�(�g��5$�4Ɣٓ�=?��j�Q�IX_�QXkEFR��
>����_�� �'�E]��dGG�о�4.IDK����u$�n�ݨ>�P
<>A;5��ŵ6��s�uc%uv��ӹ;	CO#�:3>ג����8D��SpA��Y�/zs�[�����g�Obs���^JQ'X�Z�a~���׆�${�9��I����t��~�)�Ү�U�}@��9�=�����#��.P���J��n��[�%�Y�X��A�S������n�9O)�-��M�.��!W<.�3,/�1��J�����W��lX��Y�E�ӝ�W��۔�!�Ů�ئ����\%N������(�5��b���a�v����,2�������ۚG_cr���x����Z�.z�l�|����/H,
^��v�p����S���-j�:/RU�,�=oZK��~���ِY?lYr�qkh��F�f�����Ĥj����ũ�ޗ��"UY	�ªB�=�#i���w#	��h�;#	��=I�ʑ��ٕ%����C�ܩ_�OgCR��'�/�����s�w
#�^&q�6P| ?!� ?>`���(��~��u�+���I�ٌ���i���N�ǚo�?38�B���Crw�E���kd�F8 $���2�X�މ-�ED���$=��2���Ņ��{`A��o�R�T�醧>�(KP��Ed��e��<�L6]Oa�du1Pf<�6
N��}FXov>F8E��q�o0Z5إ��bJ\-�	�W���l�큔�}�c��� P}�Ӽ@��	��Wx�� _L����M~�gD�#z���-ټvr�fS�3W��f!�A�?���6���{>~�WQ�ٿ"��)������������� ���w���^���g��%A==�K,¿v��[3��d�l�H=(�6C��\D�އ��Q�OB���{�/p���(ځh*M�CH,�`�!��|
s O�f�o�5:���o�����m��6?"��R/��ظb���|��a\c�N<�~ac�EK ��N{��6��'���5]��7
� ^�T��{�ucE�#=ǶEF{�k�$���3EF����[��K?�;��v�cՋ�xtW���G²����B�a�r�����:��Y�F)���W�G35?n�
»�s��*K,Lz����b����`~�О0�nHBJ��9$.-���y���A���R.��k�'5Yg��B!c����ױb<�8pS�6zM���U"��bh1���N�-ܿ��vG�3������w��*���an���� ����J�!�R>tB�	��nm��s�����
�E,l	ƪv�qCϵޚ6�l�x{ַC7���i���w�j3/�0�Ԣm�V��x��L�Bø]��h�3���%��@`�P%�M�D���6	��A^m��Tl�ؕ� 9$3:��y+�d�쇔_MM���_�7]��&�e�6	�	��G����_�K��6X#���1�P��b��3��e����}�p�#������7@z�:�RƵ��4� sֵ�:���AX�[D��NS֗���V��VϤ�A�#�S��c��p���s��۲QU���B�0�U5�lZ�˅����jy��Xb[�@���ye7{e'�퀞�Ѷ֚���4�w���y�u�Lô�'>�n�0���*@���U� >߬��;�un�&�N�.����P���("�.���2���-�Q�s���xoG�s���݂��f�v�:3�V;�&���qى�z�6�S�Y�ˁ��A��&WatD�r4 �����)��C1���~��g (su	3v#+P�4�`2�CfJ�����H&FO�r2�+��,�����Tu�&�׭%~$��/�}�����iEx, �{J�>���Z#���#6�Ц�.�����P��c:|`yE�ʺ<���n��h4	��|j
U[����#��&+�E"���߁��tlv(�J�_�%Q����K� �/8(X��ٍFo�`��[��[	c1D���|p�濕������$��^UDq�@�h�żM�ܩĆҖ^�R�M�5A4cu�"��i���o�G�E������i6̥�����ɾu��wE�.�C��u�/��}�]>13
�����I�?�����z�S���ꖆ�Y�3ڦ��z����Js�[���`�)D��z~w�L �x��g��|.�����T�����6�2��Ϧs����HЭ�d����k��[e��bEf�'��;���������`@��2Ы��H�B���$��o�KaSK�������3���{�@�!����<;�&�>���:[�GK ۂ��.���
�� >wNۚ��I�oo+񎀮C���c�T`?06Ih�+�~�Щ��A�T��)���aEəPO�j7�&��m�B��e����3��f��q�?�� x�[aZ�%l�Տ�����F���0��1����"i�b�(����"��[R�3c��?q�K;��D����Y����:���e�y�T��k�����J$|V?�A*�`�_��TX%��5����>���sy.��678�K��`�z�SZ� $�j4{T5q��j4����pΊ� �Ei�ut$�$k�)��5�L��ymZ�j�e>K�	�d}U��s��d������e`��J4WH���s�iƥ� 5�د,,7lC�����?NN�c=\;�	�|�n��G�
�
�2��-�Q����q�@U��H��U71d�v����$�qB^��ü��4�N>'a�[��Ѭ�S�
�K��v���4q��V�}�������B ����J{�ڕF��h���|�/�*�&�;���h�L�\���m[nl��yY��Y!G0D�a���Jc�H�z>RE�c@�D�&��h��߫�C�׮8��zJX�I�j�(�P�@*L���\/b��7z�_�j�~�:6�#�����i7�ϣ	�WJט�q�%�bNT'��_��'(��>��b�Cx�NO��>]���橶F5d#�l��!+�Y#��=�ǝ91��r��/$ZlL�Z�;Z���ˣ�����%��K�v�&��@�P�������V厌x΢M�{�{K8|RZ�3�x8����J���/!j���h"��n�-�
����!W���������7��ajB�bQYO���γ��DCK��s��®���h2���d��������Z�)g��4�{lT��>�X���Y�ΰܷ�+�z���[�<����>��(��3ߘ��S�}c7�ܝ�vD���F;[_��rvM�C���wi�7������y qe�7�#��t<^�
T�)I ��4�@#�_V�8�~F-&�Nr����
�R��R1�9��]	X��+��|&������%d������[��}s~`���K�6����W���Φ����WL�^�@z�	�~x�Ϗ�e�c�HYS�?K�24��&����竸b��s��[�<z�����O�}��,�5�j�c�����Cǒ�%p�8�Z3`	���*�k7���*���i.{�>+l�t��'g���
﹊뺍���&�92(똔J_�W�K=i�|�h��Û6��[�<��KI�Ⱥ����/!���?/�pٵ��o����A?���l	7//���!�W�%>S���V$�tFC��|�<k���d��o,J�����^*��IC�"�mL������h��K���:��'A��V��+�D�_o��Cڕa���� ~^��Jpa�Z���z7Y�4x1��l	��$`cml�Vބ��(�����n!��u�~����
���b|ߑ���h�	"���s"��j买b%�`�U�BrZÝ����`�kh7)P��n!��&��^��l��t�є�ʹ+er�����
Lrf�>3�"��z���^���`�=��Xv-����D�Y�0|{�Aw�PI,-i=S��Z�pt�g%�)��/6��r_v����1�9��K[8��'g�Y}�&��h4�5h�F���{��EU|����,��츜�ooW����=�d� ���'PBOL�#�ו?,��N�{��65�Q,�zг�"�;9�B�"�o/Y(��q�ފ��L�����]�}�e�D4 ���H|/6�ٕ����-c%��}����
4ݣ��~��e�2�����~c�tҍ�{�e��?�L�:��7Qr��)5�Z���$��j�D�\ '�yW�z���%OTIm�bئa4�o�(�����)v��~N��o�^�NË�j�ëFU�ٿ1�����g��;�3�����f�'^�mŁ,��3i�)g��{�3uԃ�-���0��*�0�O��� dK�=G�W)  �t��٠���ԥ�,|�#Ͷ��	o��:��> N�WJ؏f�b��FDP B�=����픮�G� �A���EG��s���j����6��(߭���!%�����_wW�d#�ֱk͒�Qb�f5%�ؚg�EE�q��^���w���ؿ����bfN:Q���"	���NA��t�[-�2M��r )��/��8�ʖ4I��{���f�7��b��:���t�S²� ��G��K�RKZ��Wz+?�M}�Uj���~e�Ւ�ֺJ����}��hM��zM)-tŀ=P1�}�����E�k�MҾ�U
�	��	o*I��I���m����OG����
h~ׇ�<�3�i�M�K��D"���;0���Tb�� 5��d��v��B(Ȇ�u���@5��^��V�;~^2�K�0���[��X�R�S�^�4�T4��b�h�F&�G����7� O�繒�\=ڣ���?҂VQP�a�h�b�r��^�Q�a66�B�W�z����c��(ْ�`8> 
�u�;��4��P���T��yURWO_2�Md�|��J}(�\��64����� w-��Z��S�
G�܏���2AEE ��:�ګ)�uiƬ��L�����)-ɽ���]�qy'l}*��~�eţ_c���..o�x0�*�6	��)޹h����:�}U�$RQf���[!W-8f����bl#��FV��W�t�@T�4H��Vb����)���6т�W잝����z�^��}:F�3���ǘ��A��B4�����
�����7N����q�Ɵ4Q���ϜR��i8�-6+�E�̚�j'Nߺ������㪚l}lx�a�iK�N����W�)=��V���������uz�䶫gW~����ֽ��z0��Fa��e��?��)�~�w,ZP�n�z	:T���%O�d���?W���l��aW�2C�HQ�%3+g���_��m��{Y,��#�ї?�2���o��S�k�!nS0 ԫZB�����v� �1}�Q��u��Wh���A���+�m
�v�CC2�R��!�⁬�i"4�O(��|����8�E
�gZ{�}�\��#��A�i�����;�)Z؄ H�S��bI��h�w|����3X�iY��s�T	۶�:٦[Κ\��s�(�B��(LX�ˇ%��fH	�$9�%��2���H��|_��e#�����Z,L*U��L�r��`a�EMr�ۘ�,��@eJ� d$3{%�R��ϙq$ih|�$�ZP�(�䅊��?#G��ғ�*#6*�qAb�]�X�Y ��U7x��Q��%lQ�^�m����v-��<����VĂ�b�?	��Oi(�^F�Z�|
����2�2�,��J7͟�2;E��%Y�ب��#!A^�L!ԐZ��$�j�Ś��b6G���>ܻq%
c5r*�0&R��`k~J?�I��ե�GvA�C69[�"�+�1�I)A�~0�%[΁��U���~�p`�y�_2r�@0�����O����J���ØhN�>�O@�U#>��1n��ڊ8S�7��#
�S�Yy ��� .�}�ߞ�����~u#I�y�a��DP�R����I�SOo2�4�v�6�����d%���7�%��dh�L�N��8������vz-F���{�b|i�I�� {pP��r��s�喦?��R�����e��)��bw��I�(�Or �v�dj��an` �^���K��#M�N���R���1e��W�K]8���C��}��H��Y�Yi�2ݦf�Қ�����˙H,�O}\�@� �wx���s��N��	c������G�v� K�ل��6^c���✠��#}c
��g�����ʔ}L�o��ӌ�xT�n=�����1G��BD'�ՂI�����4���^�b����b���Nhm�H=���?Vv�Z�m��J(�jd��߇�'�:t+WP?nY�[��oL���L�w<�+񑿆�,8Z�r�ã�ʛ.>�9È{������u\�ĥ3��e�A�������Ӻ�g��r`���T��O�d�%Z��&�ǫ�᤿ћ�;����튐q�Cr����Թ*t�� �s�N,rCFz�P%{���"���@��������>!��DCr"l@�~<)=���1�����>?qO�Э���5Wш��kBz�J�n�x}����M�.��|.N����ށ+�\�ǮP�� �l������B�߉Y�l���G)�s�B�B�'9Xc�K����Q�m�����J.�@�49�w��$�t�i�c�?�L2�����>5�-��~��mi|���_]�`!f��n��`�3ݪ�;CB1���)�������3&N2[KךU�9�
)`n�U���k Z�k~�턘;��h�q����^hE_ l੶f���%:3�����"��n�t�*]ˁ	b�p���z������!�Ԥq��I�f���5f���N<d
�>
���	�,1X���ؒ�V+�L��m/J��΀���Pa��Ts:e3��(��<�@�O�دa����Qu�l��c�#@�s楟����r*�#� 2����t�F:�EQaL�� .S�y�fw���������Zܥ�_�[�`|)���.?���3�0��ˡF��������w7��I��JDF���?�WO��t�,��,�q�T�Y��T�n����?��fs����p������@"~%�d�5
U7�wL�"O���1dm7sDd����i�A�%��"��Q�Oj�x�"���!�D}%��������kY��Hg�H2aO xC*Tc��|c3 ���R9��O��X�hv�
u�P��z��j��$��Z�~� �}(�G'}i%��B%j� q�Y-��Z��AN�v>��!��p��$èZ� ������@ B6����8o��. 뎂Ȭ��)� ��>~�nI���j�O��˦��"�XU��S��}rj�� ����o<*H��Gw~�0��6)*;���v�o�gK����Z��WIF���O�=�QA^�ˬ{��/��z��3!���xK���L*cy�>�/�*�<��	�p���g�g�Aq�[����'�~q��������-����˔���9t_di�ej�s鷇uƓ�^�39�p������
{���]���w-��bkg�� d�V	GW�0��:��jfp�L�9��L��<F����f���4�����0�@�����3�*�%�'hq5(u�����3��6�y��!:x�9t��m��/�EQKc�1;̍�HRJ�Ղ申--�N1P�Ŵ���횁��P��F&�\�A­��Gj��,�m��7+
u_:�&�����~�B��Ɯ�P=���!�T{��G.��z`�ր����Hm֛}w�s ⋈����B�Wą���M��p���']0clI<�2`�Z�#M�[76Ԑ�G����`,������
�/-�^�G���"���m���Ձ���>B<�_P�qr<F������8�\�[�猽�훁kO��P�bJ[A��J�/�L{�,�d�x�ʱN����}qWi����ʝ��h��(�@�_��vtM�+{TY�
Q��2ӝ����
i[>�P�M4�M8��/�^Ua�	[������s@h $�1�HP�yEc͛G唈20	�x���ds�]>̧�L��.c�~�S���4�����X��ZNţR��'WN���N��K�J�s�-,��J��i<|������Y&���R�ϻy�"\��5��-���7�Yc�W��M��I�D:`y�&�0�9���>�pwsz�U��$��.U���:U~.<-=L��I����JT��@�����f�b[��ƭ�@s�ݸ~j X�n> 	�w�l��UA�
�a��,�S���_�]ܘ�e9�>b��oHU�$�`�ɾ�/�bY�����&�VG
81�����땞��F1�8;"�1��r�!3�ޭ��5%dY�~#���k~,
MT���|=�[+F���K�-35g�I�Is�TF�b��Ȉ`�kdBa����]�-�ua(?�K�,�]ٰB�g�%t�U�����0���
 ��1c�CI�a$������u��J��Դ�ME"�5���v��c��l#^{N�, �AO#����#��8K�(���ɬ%�?��yM��Td��6��Z���C�n����#��յo����z�a��!K�!���t����!d�U-6�Ί�J�X+�P	 YX�K@�!�^�Z��q *F�4�e-c�ҙ�X�L�fO9�:�
��݀�-dI��gc�5�/��y�i<W��.bpθS�Vc�0����"���g ���$>=#�)%�AԱ�H����7�Wo�q\����q����N{����q�UݾPӉ�X�E^D*}=U|��f���σ.��N������.�N1[ � �	P
.	*`��9/nkC]�o�;Rt�vas�Tǜ�b��3�ZO5.�j�=}�g�C��3\�����	���?���F���"���:��7E�~��� \Uy�>��lB�5�Z�˃s�q�U�ʪ6Rx!B�v�$2�]>�!]�B���9j9���aL1'�*�;2�f��a*��?�ϋ@E �� c��^�/e�C=x�-2�"y�1�N���jyN:���M�G5�6���?�̰�,,���[�,�W��h6E
W-��E���4���<�Y�أ[������,�V1�j� ��4.�L"�Kе��j�Sn��b�j4ezT9��'?4��sn�b�v'������&Yh�7�S'Ț�Ԫ
�HA*���I�i"*������t$Z��@��ì��Z�[ o�偶P�0v}��S� �O�Yȕir��S�"h��Ԓ��Z0���Hߩ�,/{�'���c��L����c9��X�	��S��5+9��5�"���u.��Ŀ�Ĭ��E	�dB�����ʾ��B�����c��_%��B���mM���ȃ��\`�����c�%#;�E[d??!�
5�<�yS## ��64�Cc�|���D��׏����
Y�z����c�A�|���/�T�y�@<��O$+W.�`��~�	�2Xj���u���2h�\gq�T{��v��,<y杶�J�Z�Z/�3(!E�⦙�)6k4�����_�y�J�Ua�m��<��r I�.�c����jw  z�e\��]֏Gt\yS9�o�DtEN���m�H�-����)��b*�u�,ym5���˶��h�l�"��1|Ҕ�f䪡)�ٶ.��9-��}kF����J2�>�ό�\M0���u/���%w8E��Q�P\�A$�����h/w�9�A��_?z$$ڨ4;�a]��Z'�Y�w;a��Y�	��x�x��	B�v3�I_�y�\�I� �:�F��-�Iԉ�������.o������׀�+{������i�'�Z�Dz�Z{��?t��:݌6��R����<�+1��\�b���-��e/aq�w>�����������d�XU�&��^�u���4��K��͌�j꿫��.�;�f� ��'����6��?W�[�W�� c��$��S�h����\���J�� �m�p��t_��~���"F*W䉻eO����|�a��kz����,��x�7�p4nLv���L��Lhl��2q���mK�B?��]�W������zޞ�+��Ko��|����#j��h�I��E>�e7u��%ׁ��ˌ��D��;P�]�Fd[h���/a�s����Ha�Ƙ�1�ܧ��c�V�h��f���X��&�A�R���d���yu�9!��6>�+�']]�j�p�T"�E��K�������t[J�@�/A��S��y�$/������̫ه0�?��_����{�{��O���؟cAn&Śx�94%�{\�����t��^�ɺ(܉���D�7UV���-��h�xkϜ��xP�Hm���Rħ@{E]���>�PT|����l�r��s�G�,n��}��EI�/�b;rw6/{yWy���+=D
���.S#�����~�9���FY�� 
���P��G�B�������ۥ4�I���mE�xu�(
"0:�nd4��Lr0�Qy��5A��2�<��d��TT��|_��_P�<@����C]���7�g�?���o��}���8T��C�0���%#yS��C�G���R���h9Q���<�5f�A���� ��;Ua�^Rѧ�GS$W��!�^X�k�>�s9�����������\'Dǁ��[5����ŝhL�C<S�,���K�g�o��.ST��U�q�^����Љ3�(����1�	�b�^�ɸ�Z��U-����� Y(^����k��`F`��W�A�?�ʂ�Bj#K���E�h���L>h^X�Za��ʞ	���>5����y�(� ��dQ��=���'��=]�V��;�0��.�$��N8B��tƝ�H����UR�� p}�i&�5�G�ŝ��<[���ݩ,缮eC��^U;�\���,b�| Mq��{0�[������ISo(%<T�űX00���BU�2���^欻W�7E����U'���\Z�u���f[��(BCf��C��_�\��P�D*��!�!5".�/��R���J�d'm?��GN�,�[��U�|*9��R�F��;�� ���Qt�ڦ y�	�`^\��.�C�WX�c��##~M4����E�.�: �=�Pz1�!�ULw)r���h�s��&��ߏ���`MLW+7>jb���z+2;���y<�S���S��s�g�����Y���WTyf�`��o���))hر�~3�Eb?&|$���o}���4��(�	�12ڃ��9�uн��hz_�lE�V�D4"� R�����\��ـq��۫I�c)n�P�ڗ�r$�F�|����?UH~��E�կ���R��o_B�o����� �G��]U�\�Zi�?���gI)�ya|����D^�n��4_���n"���=�+I���q�޵��=�{P�7�/�*�a>㛤���[:S���D�ה��`��bT��ic߉��K�.���I3�q�9z�\���ܖ��苔E�G���Q���j[hg��_���37����t�������lĀV�DOK��w'�:Ɛ��2��,�*��[����>Y����E<i:}7���!��!,��x�y��.>]c�E�/s8e�^���r�Qc���&5���G��&���U��\��\HL����bp>�	��\y�&ZVs�`{y��m4':.`�L�u|x�[�y��x����©��� g���[mz��e��S�|({`/�3�Մۣ�-����1u�ß����`�9��6C�K��FR����+���$��z��Mz3Ʋhv����|7H������f>d��:�U�)�ڬ���ڂ���b4�� h w���t���%hsKsٖ;�B�A���2�G���g*�w���y�V�#���3Q{^���@+�c�x���^`��$\-V�/7���*�B$��])�e?���ߛwlWt?��
�ɠ�{�^�^�yO�vwe�����+Pnkzb笺us]�>^+ߜ�̹��#H���$�����?��n�i�Fm<+�C��u���O��c@�X���ku/����1ÝPx��/6r/�HI��PV|MZv��n�ة���9dȤr84���]���wM�@�D����5�Z��F_�6�C"SH�4� ���ǥ�!-��u���T7��E{n�۬�G�(�b X�ڋ����P��������zC�6�'d�ۄO#ך�~��J�Qo+?\
#e��qu�޻�p�G��4r�9��7[�S��w�F#�̄�o��mg�
�2��9��b�L�/Ê"ޢP���b���H́i��fk5����w�9x�v�X�`�$� �a�����.5|�a|JKx�}��vfLI܇7T/�
N�'�;�k���x��.n�C+*m��0�UMQ�j�*��b�dD���ޕ�r�����c쐙l��u�Ox�g�Y��L�U�k��)(!)8@�}�X
N-�~����7��`�h<�׍��4Vj��,c/򎢍�!&K^\�������Ô��ֶ~�\v��B�o�r�h�F��L~t�o<B�3%K�!���ӗ^�HTD��{�dY£(7ā��(����K��Q��=G��ٔ�Qؾ,J��C�
��F�����<��9*S[-��QiiD@�����_�ډ���W�	�ڼQ�;�U�X��쐆"����	%�g03��"��W��\U|/���v�+-k��}����0cG�;�y��]9;�22苣������+�e���'�2�B�9q ��ȧ���QL� k_����V>l��	�sUؕ%D����1�m:�g������m��|q�º�S�������t/M'\z�ZL|+��������o#?�ɛoay�IŮnۄEJGT�2�d3�h���}O����*��Y�u�mI���=@�螸�rjL���|L���Ť�"%�ϝ{M��S�RJ�x:��c�<�77!��X���?f�SR�i���U�/)�˫UǶ�;�({�4��!9V
���]ԋЃ��Ɍ������[�I/
ڦ.�ӯx�~ݹF/�Ğ�S���I9S�}��	�4����S]�ձ�&�B`�0����V�r|�f�0���21S�B�����`�Ϲ�I��V����Þ[����-/ǽ-:M���.�x���{�؇���H��Vr�� ��H�OyѼxĄ%���c�	G����@�v�LИ|���.X��D[�'�U��x]�����LՕc��$C��|�Q�ai���=NTi�ϟ�[~�z����ԝG�$���֕�(�W|�r�΢��n�gp�qQj/<��]�)��f���E��H�) Vkދ����/^�&��ˣX�;U���mgΌ�Z}FD�K�7�����R��4nţ	�|r穁yaT��qpɌ�ߒ�Tfz���h��ǲ�� �c�4R\��T��&�@�;B~gU&6���W�8V�\�w��U`o^B�S}�ޜ�r�ט��G���||�U��0�R��{�N�)1�:~b8�'ә�I�ğ�j����Â�E��a�/��L��sm�Md�kH���B�������t���������c$�U'�r��e,+~V[��P�t�#}�Q�c��[�y�� _�4�y�����5���B\��z�P���ܔ��%̴º�8�o"�%d�rzɾ�-́ak��_h]k�1�!H�D�[E��3ú�D8�v��fq����je���YJH=�i*:��|u�2��������[:v�`V��Ѱ��yUD�<sq�����%t8��ڇw�`��$F����2=)��G�$���d��@؇� z^���0���c"���l��㗢9�pI��&Zl�m���H�6վ����x��{.��]��K��a*�qN���>�#�AX�>g��� ��)��"hȉ��,+��(`�7�c�QL��Ă2�Ӣ�UO]@� Zj��zM���<s}�A[�JL�ҮzY�ƀ��6{�\���Jԅ�n��\���1Z}�u#�p�߀�k�m�gϦ*A�o����k����NL���(TH�x��m���
��[_�o�F��p���8�`�kI��*�R�a��M�X��
�Vu��l�A,���w�~��6W��:t�Sp
�Z|���Y��M��39T��M3H�w"�V0}~1v���BarQ1������B�3_��?�X�D�I�w���ݦ�t������П���Ƙ3����Z�;me������1ieb"��"V�r�2����7:���oYb��~��|����	�F7���p�|�L1�{(��7�[gF���N��%�v�<}͞��u�;T�G�U�A#�+�}i��,���?QC�p%����|zҜZ��ղ;�
 ��iîo��Wה��3m �((5��z��~�}���X��\�'���5sKu{��Nd��-����9���!Nt�=VE@�h�"$�������X�Iƥ��a~��3~���<9+yׂR��3�c�O�MV|�-��ߡ�~��U�RZJ�{*/q��'%��z��I@�o�
�2�$�{�]O����0Q���:�=���K;e�tl�Ba�����-�H��I�R�'��mq>Ճ3 �|��
q�,n�a�hE!Fs�r����Ko�d�Y�H�[�C�w"9�<:Բ�5h9;,;�D��� ���^ܧ�"b¼�sbR=Rf�mF�)�"{rd�JZdZ�e-A�ݏ�0���p�YI&�Lt���giɦ��c��E��C�h�=>���.1r�i���KW�4.J�k怹��(v8Y�!QU��&H��K���_e$�+؎�YѴ:q��Z��>����AW"ܺ�·������K�L����o�e����?��ru�".8"'��4_�,��kz���rg����s"Oy=#�;M`�4/�*��B11B����}�"���	�?���]��X�)=Ñ��pֺ�Ǧ�G���4b�P�6G<��*!r�\O&#�m<b��3TL�D.���$8�����%�"�|+�rH���Ş���!���P��v��ٝ�!A���iN�]u[��q�[��mT����74��H?:)�5�pp�#�e(��\��h� ����zY{W���=��T�Z뉕U�@ ]䠇�鼠j�=x��1MlCd�O��^��O1�923��h&�p�S$�/0[:�Ҩ}6�a��y=gU\��5q�o��F�!G*�Y�����C�]_����_����V���W;� ĝ4���V)�i$��6�G��{F�O�J��ޱ��nf�� ���>=x��~�z`^�*�78'�KVf�@�X&F�l�`v?��.���������˅�����g��(�.T ����	�'q��ox��v��V4�R�'X�Y�N�����;��/���2<(�=ϲ�C�E�O����Ǭ�08�ه�p�K����D���u�9U갹�R �)��%�̄����a%�s�.X`㥌$�jmd�_w#V}�U��ˤˁ�^F`��&�?W���Y�������*c�� ���V;��R�ӯ'��|��r���\m�P}WNj{/8�1�
����N�(ԠN&{kgK�2*	䀆� �ܙ��s����N���Q;_�'��0�t\�R�,��n�DE,�}�;L�7y�e�:o�x���bj�3�W�K3�1���_ �Uͼ�q����L��,��^�/��xWy�����P�<-Z�ht��f�PI؊���36�q+э�?�VCUe��Px�d�K|�`����g�� B�1����1;H޼���@��{oe�\����Z�O�}e��\yHoړz��)�b�5�����E�7�x��;:�Y��ߧ��T.���� ���*�4T9��1��&e��2T����V��M3�J��\���}fD+J�M����]i�����̝
���<B �rJ��K��m�ϽW������:�C���g����Aد_n�� ¢�7G�{�Q�0�n��,���nS����
�$Ý�#��P[$)I9�p[M�������)���7�W���bF_�`73��Re�{�;�ٵ�����\���Ny���Et����*
v� ��%�����4̚5����ҧ�}�{�?=�^�J�ʌh������Nuk��s�s��r��h/��7$�8F��8
5v4@_ZE峛<�cy����aX>��4������&�5�e�%2+��?{���Z]�_�D�YN�ĸl0�W�H6�	����*�����-	��h��Q�1	�R�R~F)ؔ����nk�9I����N�{Qrn._����D�ڧ��ۺ4�-Z!�o
w� � �c�\���$����>,8+���Ӡj�w,]�++B��y.����G9�S�
30�ww��K̑�o�6�-�2U�[���J0�o����՟���l��#kߩ�e��|��n3�I�y�]��K�Jg���#�;Q���^�ώ%xJ[��p�%���=ޚ��G���JJ�2�g����{��}1/<�ԁם?H�l�S���>�^JU=AP�����@��pR-^]U���k��E��K{!_�?:�13���`���V"kZ�خ\	��^��ʇ�m?lX�Iњ�}�W��3��v��%'�۰v �Mz^X����=�e�E��������G.���c�-��Bm�Q��c-�im�V2pߌ���\
J��u����KnK20��*����J%>a����%�Cl��Ι�A��hg6Ff�k쏐��*?z��|���;��0�\���=5����B�a�
���þ$���L��O;��~�7"����Mk��9�:��uj�W)ܴ�՟�fa�� a��"�5��';s�{~�~A\x��G�Y�W&~�f�/=Q	�c�)G��a�z� s���a�c�m(������G�疋�
��6�C������Ow���s�� ��b�6t!���y-��cO�K,��R�`���qo�h2��?�C�`���#�'f�~iD?��D�R@9�5�ຶ�^'�l��͖��._L U?2X��d��w��,��A��<s}��4y4!�t�J��TO�"ήV�0$6s���8�X���X3d���pЙם���2].ռ�H���>x�����~�5����/-���$�ڥ�CB}�k��͔C����t�~��6f=��/��p{o��3I0Xk	�
@�E��m-Q����?�����j6Q���i:�?�����lcg@McZå�0]��#�r܈ho��X�W��Ұ��ǅ�ru6w&k�n@	�
�֊-D�����t�Q�s?��[��S����W��cI*�	�z�!�$�����z��v̬O[̫�W�9e�@�o`�n���o�8������mgk��5����&ݍ��l]?p9+]w���0� W�Ɖ�h6�D��YpT[�9<s)�����Mdl�ڣpٳˀ��q���O��aZ*x��}�.E�ޔg&��G�뻄���P+F�+kl�T[۱O�.q�l"��s�׍�KR�Z�C�F���1�jnS����}��(bl���@�3��k�2K�� i25�/;ߑ�?;����� ���ǅ&`I�"[����'
^�@*z�и���m�s_����,fnGS��&&�nl�����2\�ۭ�r��0w	��I�q� ���cJz�����U�Ħ���0[n v��u&2�"�����Cڨ8�D��=l�t(��u��łh��:�9R�pn;Lͨ&��Ƌ[��M�#�$Y]�&�<����`{&�<�К��JRY�&r�j0�Ԇ/����c���ͨ��p�ÍrR/��ke4<����\��ѯX��ȵZ{ t�N܀@�\Lȡ�p,n��1��f �#f�};ܲ��̓n���y�����������[ұ6 �54�e�` �԰=���s�!sB�N͊��B;ք7AH@��k(�!�?dx��v��ئB��tf�zm��4M��Cz�mRKA�F�C�'ԛ9W��Ӏk��i�5�Y�ĳM{6(�2�8Q~+�L��n�����-ᔪ�R?S{2�v~��&XJV��p�F�-� ���->٫U�0�5�����l��0���~��!J�Oۢ&hŞWr�%�NA]P]�0�h8H�e�1����>B�"\j���f�f��şuv1[���Ο-T(η������vQ�c.��o�����R�-�-v-�.힩�`�Dx��lZ ���/j�v!�/�ᑼǏh��ҥ�-�J4� < ���3����7�_�~�.�j�wٿ���o��0��/Լ�����*fC��.J��"��+F�v�|���O�ig���v�����7mtd��[>�j��nDpP�"�<�b�N��uJ�/ʅ�!��>��K��65A��	8�-i*�K|���
���6^�>���m�ifQ<]L���)�d����WJ�gQ���T@�3��1�H���+����<~�fh�x�6~T�^N15{��Tw�#p �(-�[��;�VZYb�iD�p@A�<{��h|���7#
r���st���9<eo�������E��@u3m~Mݗ<�0���3�O����3ب�?��-�G��M!�z�t,�_�w�)� ��ۙ�T��{>�=?��%|%��<���4����FP�B�0D���!�'�m���uYD~�¶<Y���ig/go�ˀ�b&�-�
HY'+�������jm.�����\cj[;9c,͋�>>&r�0����~��q��o*Ш��A�v"�MECȳ�Z���8���� ��U�K���eɯk����~�&,���l�#jE������"޼pu��37 N���O�ş���{�����iU��Z�t� �S׿�XK��M|b��J�;cK+�D���;���Afg����`�]T�kA�$RW<h�O
�Xi��C��G3��{��0�1��*����ux�O^"�Q����/���E1��OS5��	�G���F�y� M3xy��-?ʏRD۵�����s���J)�R׉Y�	��7��0ANu?� ޒ�b��c��oש��.F��%=���c�u�K_جσ��~/w�Xa bԠ�+�K�
'�)ħ~žؼ��8LM��ID��K�7�`w\�,�Z�U;�P�MKܾ�I��>��5X=�/�!i1���5h����s�R�������<!�,oJNK��Ҏ�@Dak�shu&�[f��y��ny��>�R��[Ӹ�{bun��\㴽��3��F��o<%�
��soi��[~�����0?-9��q5���+fU��G�"�ꐨg7�,Ҹ�_����U6}�Sۻ�������z�cC�/`[U�^T=o=uЂ�ў}�'�B��L�ψD0N8h$�!;d�?c��4�z�y�g������a|��r����B]1P�o���@W��ܝ���B��������If"�y�*���+�q_2��+��e�A
����p�{�F�4��!��.#;ob�zv�6�>A6J	J�A�NUWǗ:tr�n�ZĴ��P+6��|��Z��)V�h\,h4��aj\!�6�P�j��f�D9��q9��Þ�����t2U �y�B�<baƀZZ�,2F(L���y����Nk0���H͆_T��%��3�����; ��M$"7�W.L�3��먇��ܤ��m�y5] ��N���	�i����[r��F~}�8�W�I�?�y"sX��j,T/��G���n��A^���j��`��:v8l>��9�(�[��H�0S�h'�81�������g�6��^O� �qc�" ��'�F*"�����������+a>��n��็6[g�8����i�6����(�K\{�c6W�<��8��>�x��[�Qޠ�n�Y�� ��U,he�Rs(�L@�ŋO}�Pnl|`9E3k*��3:�E�jo�_q	W)Զ{��A]���q�����l�R�6�鱨G�bmԦ��%��' �Ǎ_�Zi˼=�Ţ	L{q�y6Ƴ��u"�ў��W�ͳ2��~A��qK�����NYu:���ҪuJQ3�Jn|] Ӭ�� ��q��ϓ��`��W5T�"V�kp�'��f������