��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��,�y�}�ǰ�=4d�H���`I"��W�`r���T:tB�T4D�m�)�	1��I�t��
��8(�8t>s)ו�."[�漆���]�~�]��;�O(1#5�-� 偙O��QZ��~rL'�x[�i,mׇp���O�I43��4d�,�H�����SN��d���3���r��m���̨T�I;uj2Y� Er�*p�Q$Gm���p�V�`�2^���,hz�<p��l�Bxt�5��s��\yq���#�@W���f:m��T�	,*�񞭋����_��㧋l�	�\�:��uGd��PǷ��N�I��_����Tuv� ���us�(H�~�{2H�:Zor�Q	#%�3ˠ!��iS��95�,?�.���/�F�i{#���Tp5����Ҥ0{%���2vpn���X�����@l����3dc�ק�3	�Ed&3�ZN O���z��s�yxӡt��v*}ԫy nj#��lc��m戭k[��5)�A#�����8�!�]�Z�s�M���t��w�!��'ÒE�rv��Ϝ�c@<U��\tq+��&|�&X1)C�����r�A~��B�&�����s�:n{p��͠R�X⺂L^��R����c���f��J^?��ܣR�O 1�rV���:��T�4���AD����˩�F�w��)Dm�O�b,�a���1$��c��7t[i2>�ޔ0,S���󧇳Ϟ�ᒨ�-��}�!6��Jyv�醊�^_�(�H�(y^����o#����X��3-�k\8�M�T�"`R�DF6ȕ� �,5�;Ҭ C�k���1\������k�t־9�}���� ���QHF��"��t�9 ?��{E_�7��!����](�S��0�q��w�9��=�i]�1�GʦȪc�W�XC�|�$��}q�6����zf(����լml�dz������*�eLD�*�,�m�]ہ6����D�Gw� �g��' A��)�m���b��ӎ���o�6ūvO��=�W�������}��	����z
��z�&�P�K#�^Qץ�_������&�)�ٺ���/��U���WX�wK³��4�d{B9/��&�	�d �Y ����6��-�X��o0O6K�-آ6�F�,H+B�*�5	��~��6�q�?T8F��Ýt��_Kf��b�Myz}���%�l���)�|��za�ӗ*���>Tk��EU�[��2�Lu�uU��=��L��Vn����$a�9�f~U=w��h�l��r�7eg�1���$��=?	)�Q��^��(�OɦǤѲu����u�r\QD��q��ɂ{P��{��d�G`j�'��fB_�R��.Om:�����Xk�Qn����*�h!�i^p)�\n���H��;?�g�x�����ؗ��3w� 3zED�ͪ��h� Hm	��0I�>�V\�V���1U��:~�Xa��P�ȴ����۹@���`�����h�s�y�Ph9�P��#� �ҋ��,Ne6��0�*����p���'z���7��.��<�A̍����[2@G�����F�'�#�����*���]|����S
B}�5�D��K�u0|��<o��)KpV�0��tB �߄8��v�x ��Rb��k��� ��b�(	���^*�\��P�t@1[�b�u�7eyV3LIlN�xP�[��oig���u���"�}��z F�i��x&M���L�1}*��u��1pP���k9N-���h������'G�JcN��ҧ����ީ�U/3jX���q�gzܞ�
����N8>�2����v��^nH���)+Ÿ��'�|b�::Z�&����r��o���l����������Zk���ܿ�%u�Y3b+]�p���a�1�)�"l;,.}d�Q���wl �6u��̨�h%W�.z�]��aN�R;D�L�L f��-5�hHJ5V�`&��<�Fc}h�/y��u��s�86
���+��iKr��Η�)٪�
��wěU�h=�o�Q�) x�ymP��)�qa
�~�$���l�s�3t��d:���k(��C���@5�
u+�4��3a�WTO��Q?�A�z�jG���&�p@D!��dbZE�@�=�#m s�k���5�ms�[�k�U�V�|��C�<A��oRu'i�܋1��J�q>i]i۽<`�,��u�FIF3R�(�A��o��r)1�wWQ������1�z�A.�CD�ۢ��Z��O]
�=�/���01c��Z��`���)���ܳ:H��O�\���J�Б^� p���L�KVַ��3HLѪt���P3�����P���2���-�_ƕ9�yG��#R*�Cd��	�y�(i܇`?g>S���t���!�`�x|>��-X��]O��9��V���c�U�"p���,���MlM霠��������O�����̯왵fyKf�2h�Pa�.�#s���-$�2�d�_E�|�a���P���j#d� :7�$�?� 9�-%�D
�Pjކn���Vb�Y���񁸿'�=��{��d�h/�^�t�Qv�7�RM�.T\fA�;ך`�U��tf��Gƍ×w���)w�M[���9r�{[�aJ:)2�AEM�琕I&�<fW�1�
l��J9�t�=Fxk9jĈ«��y�h�����xNKA�����o�bO�F�p�O�L���k��Gk��P���K��+��G�k��T�v������C�G4�*�����?��ލ�cbv��gj,@GN"\��!���w���Ո�g�>-|���'3|W��=x
���m���c��I���]A�]jA`	2f�m�I�G<�*g���'�0<�m�(9_12r�s*��Y�i��1��5zg_�����(5����7ܦ�R�h�T�����p}	��)�z�gv�?�"�m�ݩ�ι/�d��-9?W,�J�Ҕ8����}̠I|��i����r��Irg�Es�t��)�?�;����}(O�5�2(��D�Qm��0��Y��P{l�dSk�����߾��SRte�o7�ئ��ľ0$� �@6��]Su��6K�6��!B��~��N_��̘\O�����C3�]L�^i�ƒ��W��vC��C���'��0r��@u����I����K^@�[������5m�(�M�W�[�_i��Z�k��_��uG�kѡu|C��'y,�$����p�JO;;������SL���-������Fr��f/��r�R��Ʃ̰<i���BP��y��m��TJ*�E���-��s�,�yy�����O�kU�F~�� F�(� I���tq"�Xm�͵�>��J;LY!!/��h*�fǏW�%��
2�:��0s���z1�v��i�t~9��HE���n��
�f&m­����������Qi/��r(cI�w]ɰ��"4���ِ���7�1��5���t�qz;�Pj2lHV��t..=�(�ǩ���2>;z��إW��CSAt7���$�@/hJ�p�DI��T̐�1��Y��o����)���i{�g�Yl�����϶�ꕆʄ�Q51O�R�8��=G Q�6�1�u/ۨ��4�U;߁���d�JHQ��ڲ���꾑�ց>k!=���t����� #щ��Dj��kF��s��6������֭����ѳ��<�'q���(�^K��(��cy�Sa�]j��jؗO�~�	�*��K�SM!�eQx �+Ց�S��֐�x�����bnq�v��l^�^�)�� ���BxQW��f �Y'���FYP��뚡��xb�7�h;��¸S��B�br�������K��T�����������.z2�{�p�g͜kr�E�AX�X,)�����Y����._��h�é����V�j��0��_ނʬ���I�	��iݍP�)�����W9���d�P׌��9��bz��(�Ђ��6B5�_�qP�0�;��ҷ�H�� #�_!��\�����ϔ�[}�V�Mf�H�<�ml[kE����c�#�!U|���'�ry6�X���r	�Ǥ�ی+MO]��A]Vԕ�8j�'qZ�qr�{�zbd�[�l9A�~�VzS-����x���뒙�����~���=보{�l�v{��AP{��������̽#�N��3^��T;��^{� �:��K�e�d�qs�?n���\�l0�@�څ�R-��֨�D	�L�����
j��]�r��T]��w���հ��t���C�ܸ�G'N���s�W�KH<Y@N��lN�aV���h����Ԩ [v�mZ��l���@�aMk�_�h\T{��I 73�Jo���.[�[cj�K�WK��Pgy�핡�-j�q@���j����V�W}M	��Ə�jå�I�s�4f}X��2ᛉ B�"�.T�Chi��S�@;��X���Z�j���o6X�}ER������;���[��<ԹՆ��M@P�/�w?�ɵh5S���=�����ۉ�]i�$Sd���*���c�M�H`��Ĭ=�iE%����Ŧ_��w_4�[
pMnTj�
,|{�������
Yz	�d�� �:h�͒DQ1}Hv��۽6O���M��ӪA��SN���H��T�CS�hO1�o6��\��^��$NM���7[�"�z��-�#�b�r;�K�@�����HV�`RhA	g��r����R%Y"���oŎ�n�9��擁'��J1���+���ܞ5|��`z��jb�{]���!�P��i4L���~S��)�`U�a�4��.�2xXū X׶��WŦ[���6�-AĀ5�?V�_����'�>����t�k3|T,�-��CM� \�}�!��Dَ?�h�>���I/m��#C�%d|RF���FU��t9����wN�ZӔ�����|��^Ⱥ�pj��
f�m�н�YU��.�����%���#�:��C���F DPZ�]��O��� �����4��Ɯ�AU��S��.�I�l�s�>P
�%'�"��s����>��2��6A/�M����S��)���#)�;�J/��Ӻb�5�j]�]�g,ʿĥ���J�����ʋ-l;��'�j��͒cu�>ɷ��3T�EXg�8(�:H�:�����y�ړ�Og<I��#5W)Ɇ~%�,�Dڭ*i�H���_�~�QF�ȣ��z�����֩ŝ��Т�N��`{�Ɔ�)��Ӯ��XE �$�j��0�eU� �V���.XIb�iy�kA���?4��C�ߐ�'/��.w?}[���4��j�#pQ�����'vN�t3Y�Y�!::��e9�~NXdc(b��SM�'�o�������"��`�u��%�;��A��1�=☏����.���[ld�3����\;�st�	��i޲�
�H�\o�z�Lί(o��?/����̀*\�d2^У�~���[��M���.��[��9��x��F�#��G�O��J)}��&�?����+-مic���r�g��hIA�l���ៀ)p��֕J��d��' vmL�gJ�^c���G�E��M��&�� w���$��.W��FM�wM�5�(��N-,3�c�kq����]@j�����Z�5�ϳn��q���q|zz��f�R%�6=,�*7��j����
�8k&/=CC\;��`��C�<��*�
Xb�[�X15~�~39��= `������fm:/��j��R��~P!����Ȏ:�ߌۋ�� ��h���03�x�ځ�^��Ω���&^�12J�iIZ`ӄ��h+�U��[ſ>0�@�D�v�~��efWZ2\��2��3ȹ
@�%�k�	�Lpj_��1ڽY����{���\IBZ16P;"_�A�$�xH"2�GEѯ.���;�L��t��_i�\���s8AS� lO%hhub�.�;q����Z2u��Mv i�D/S�~�v���8�Uh /�uC5�}�~^�J����1�鏟[ak;.���G��q��&C>��Cq����O	XhA�$P����+fua���i���^b�'ݝ��&T�Z����}D�f�8ci�:��_I�Y���j��Dʨ�=n��y��'��Vt\	qבj��8�x�s�Mt����~k��T�AQ���W������p{�.&�E�Ǵ�S���~�#>I�B+�P�z.�E�2�.��|u���!6}��p���3�B�RvA�dt:���҃��7��!�+yW1x���^��G�#��?�D��f�������S�'�j���U�i�,v=Yt|!Z�;e��=7"�7��{�ʘ[�����m��|~rK�� ܮ󯛥h�ᷱ�� fA�H7t1-j�M]��\�U�]�-�f��8�1n)�j����!㉑��<��{@/��jr(�m�!٢�)=�����P�#-���q;��3dp�M��EŦr�q I�T��7���|P��	y��uӸ�����r>���p����4z���fK�&�͌%��t^�%��|u���B�I) {��]���H�w0_�%���N���p����r���F|u�q�@d2�0�$�0z�=�@���N0�<�#���	κ�B��X�ࠆ�V{Q�A�?���46��m��� 9�����O�;`,X�y��j��f(��S��yǊ�4�۽=�{2d�#\��.7�Ѱ�ί�B4�C �y�}���ء��Y�zz�Z��>��O�,&Yg� �h(s|>� ��~�	���؊Ѐ�*�έݯAoSDEcY�϶5qU�Ǳ�dgT�%��MZ��� ?��'<R��q�LRiE�މ�S��SX�X;Oz��9;�`ԭ��kyj�+g"4�YH�~>��aw�O�=�ZF@� ���c�R�=-�Y1�q��b-�����L��Ӧ)L� ��f�R��5�:�b���+��f��(z"Y&�����!.���V���+Z��i����a�D����oG�&�+H�W �in����[�#����M{��Y	��vT��{��i��a�y�z��вsA_�+��bf:%W�U�le��o#��C��{���J3I�C�+�&��ͼ:o�1p%TK]M�#�v���R��Q�r���_�6������a����9M)�@���(<Ϊ����NE��E�^����4�Č7?��b�|���Yt��Wc�j�ɔ��>3���gQ�#$��3� !��'�%��eO���`1�-�gW�G}�G�l.�7wxŢ[���f#�w� i�u��l�%�i��@`����?nG�clrX����5����5���ʟ$y���R>g��<˥9�������=ցB}j�=y�"m��hI�#@�}�4�$�@��>*��5�-�אw��t�fD��Τ����n�1�`X���Y�|� �L*L���� �F�CZ�zi*n��j��ņ�(�,ǳ��Ǘ�h[�Q	|�:�a��}��i(���Q�(�_��D������=�v�h��bql��.��a`���I-��3��N�>^ݷ�]��É����Ҙ�3�ю|���F|����X}����o��-I����]l�v��c�C<��vh�[0/���F�2��X��{ގ�g�ZD_#��M3��`��i����c�'����A����Dd�c��m�-G��S�qơx#Q�_]���6#�z|E^]����N.�xi5��K�Ύ{�}���4h���	d�}��ܾ��|\﫹l=36��u�]%��s8��l����c�gd獶`t��E�}��@ӓ�Q�����WN�$hwW7����Mx�=Nv�`�����}ܙ!��]�x�7�
�B��J�&�������(}�}�|�_��ڷŝ*z�ϭg���^����ZI����
�u����������.�UE���'�2U-�����V�@^D���)vUR
!c9>k$V�{�~���61@_�1�ut[�6�Oa��Io|�b#F���G�;>�X|�S�f;����'܋��hu�?`ł
>�FK��ed	�����ǲ(��/��)p"�,^l�[���cm�Ŝ%ʵ&<r� �O);M�[Gi��ƌ4:[o�E"�Go�>��{���'�j�zJS����e��#��3C��l������Fj��d�S&�+I�0��X�ƒ��\���\��tn�h1n�l��K��B�l��8���s{)W�j*�6�b��������91����T��ѓJ��j9;��I��r���Ƽ7b��E	�`�1�u��]>��|�q�z���НL���K�{�(�$a�@��൨�'�!n�#PwEŇ~|�f���7_����Q�����s�/T��u�:R[$rqT�7�bF�>��D��~<�<!�)�W\HUb
�6^G�\��T����}��Y]��9Z�hC�ໞգ��e�⁑�S��,|�pO3F��.����g7��%_���:�{w`t�Vg����s���	�����z�A+_M���Q��+W\�ʪ�@K�ђe��c _�\-�"U*��<Q�w~�o���̉�U�`Nv	���L�d�$�D��g��<�40�an4�Վu��<}`����W����gM��Y�(E���D��Y�Z�t���(j���������ju2/}�'�3�p�`I,��!��^���`���<ɐ 0Ԅ�j!�9��n��h��m�y�R?��5UBwƇ�����F�1}��@�Fʨ�/'���%��m��2|�^Γ�Ju��G����Hh����n.>��]H/������N��a,t�~A�}���y�k�}�����SM�&�NmF���R�)��5��o�@y�_��P�ۋ�U}�� &���~�K@+g�6��w��5 T����˘tHm_�k�;Goc(1_�Ѫ�j��	 ����t�4�	�28@=�B/��O(�yZ�z}�ͮ��ȂL-�|���d�-KS����wؖ[����y���.U����	��Xk��k�瘼�,�&h�v.�M�2&N1�V����LP��:p=4������E04���A���+ �'���&��
�h���9.,�d`
	?yw)�l'*�������>�`����V',*m�s��G:0q+���м9FY{���I�mh^�Bj���5�m������sR�(�A�Ƈ�{���+���C`���Pb���pt��B����T�6��y�%��_>��>��Q�r&@�a8^�@[9��"��,s9�|�+8���?�)h(⥳� �Y�[t��+�uivL1~��y� ��x�iQ]�p�$ǆ�$Rc�@#�+籙v3N�/�\����aC�K�r�Fv�vJ�:iJe.by`���%����SF H��8�M	��ZF����Ha�.�e���Y��|\��@[�b��K�8��8�P�F�B�k�Y̺��� f�.ܳx^A���rG���p�9Ǎ�^Z����+�癓�W�ʏR|�c#��gNv�]O��ؼ��-�7����q<z��N�*��,8��pC�:*�����C�-����и�b9�1����0a/ӧ]���Aw[,��=�~�#rD��:�m�8��k�Y�Aܰ�;����y煃wf��Y̑L��P�Ck�O�2Ǿ")�1ޝ<��*��S+��[���z?3L��e?�_ٍ@�$�!�g�"���yM�1�> �%�S����rF�����=2V�oL�e�<9��N����@���02I��,�p��DX��X�pV4qޚ���L}D��ms�$$[|T/�#�f.P�=��5�O�y�l�7������fsq �JJ�,:����MH�����(_'�C�y��Z&	X��V���&�U)��7��u�����`�ȱ�$�=���\��q��s��us�x��߁�.�dvɩ���~�J"�n���94xvD��'IZ9AJ���u��E�������M�;E��n8	zFdy�j���e_��]Z͌�e��`��=�~r9I����S��G�5WD�3uQ���VcRR����3��r�?�P���=	yeҷ9�>@/�hIƁ
<?��9}����X�i�hpz��Jx��[F�n����݂�;$��u��$����ӄ$�xTB��Q.Yl볥�,�"�����i� {HV	�x��Y
sq�{#7C}#����_$�����<o�F��ZE��+����$�e���
Yn��K	V�]5���($H��^�������Y5�앬YQ�t������M=�Մ�b�h�Ԣ��)�fp��T��+�����w�t�*F1����>t������^2�3�g������%E%ܸ��`V�EE}+�pF�;Ht��ܸ���3'JS؏9�����b�����bO竅�\�5�O��{����>̻���'(7E��8uu��� �(J���C�=ͫ�#�sj{(�TVa���v���vZΣA�f8#�W+R�����Ӹ,�7Sa�_���I.X�Ss;�ڝL��6a��9Jʫ%K��a�{�/�1ы'��
Q��`1��]�Px��6�1汁�(ZŷG���|�[�}��P)㪤4�rkE5��!7�v�:��A�'o��p_�����8��6:p�NmW���{���]����(�h�܈����|�M)�D����?�0	_h��mg(qBמ� f{���Wͅo��!�A%!bBiz����j<������x�.�-�ɗl�1q�RD��& w��U&��Z��~��ux"�b��$�^���[�~P�����JC��,/�Y�/�-b꺡4u@�2}��_Ƴ+� e�Sf��1�X� HRm)�VE`�#��NU�9*.>}ͫb�w*g���7(�gV]�CW*�Ǖ���h`��@���S4�T�~ >������w��g%5�j���i.��nE�7VTj�����LI�V�PM]���Nѹ��u�A�M.�_����\�'r͈ܦ�����U���3C����1f��RO�梸r�+�����kw���*�o���.��'�z��`���Q�-Nz��w��z�rh\{=���p�f��3�H��k	u�li�eOB<[FY��M]����<�ΏW�`s��$߉��w�F�E��pdoRw�����vO�f(��?*	�Ro��R<DY0��h\�`АQ�\���B=�����f2�,�������݀J5Sa��#T��3���.��V�
�Xy���N��Q��4�z~C�GP����v�X��8�T#݉y��(�� 0r������B�g�o2�3L��b/�%T6��,�����}S�ט�C<��0~���A�^�� �8/�nZ�ك�$
���Vo�`���T��i��=d5)e����Ds�����q9>�NtÅ���&D�&*��N�C����=HI�h�r��<�͔�[��m���g��ܭ�SE� �l��Z�cm�W?p"b<�5�D�;�q�ÙE��	C�Q���z�x��D�3��x��c][s���?���{r�� \�)��k����q]xe��0�(�'�JoX�#ߖsX-v���w}�MI -�~��@��.\M��|����_��-���﷒(0A\���~� ���ŕ����b�S��[J����y�T���1���abm{���L��_\k<��29_�M�P�j�2J(��C�!�R���}����pe��o��$�gM���s�=s� �T�%�1����,��C�OB3���O���\��?k��������q���ު�$�4;�J���8v?�7��]q�uy	\��e���߭r2|��U-1�J�\����^UEg|^��a��Gr�}s�
ڧfB�v9���g�3i���3���J�Ź�Ӽ!yA������B�s[n�Jyr$�R��E�0?T��{��Ujs�ҳ���$���g���c2�X ��NΟh��	V��7T��I����(���x;� ���d���� �ݙ�Y���z���k�;"�Iy�n�~^x��WY"�,�j1C�y^�3pT0��a9�L��E[��]!�8r�q;I-�{�,<�2H��³u@�I`>�}���̑� mml�vNFk�(Z�*�B�|���Je�
R����ik� nr.����������+0D"v�c��X�Y���>�)a��>�Q4\G�C@�&����?&ImF2����j�J��R�y��Ѽi��Ne���y����P�̆����A��&���-�3��݅��U�i)�K���ir����j�<��ek�qG< [�ߖ|$
@���\� �M9�3e�}#���&]�?����\�*��)��F�C*�Ҙڥmϫ{��W+�/j�n�'N\����T#���'MR%�	��gw�;�E�}�X���Y*��W�Z xtP�XSG�m/��h��shʘ$��Y�)Lm»! �Ԍ�"��Ld`�oW��f�j�N	(���ܶ�3K0��\EK٬$xK�����8�U!=�!	�cƞ�.F�d���?dY<�Ƭ�@E1{"���*���Gc�ܬ/�F��E�����K���<���3�u7f(����]��;��*��P�^�ʕ`S_�w�	��ii�Gؚ�����.PC��~B���5o�YO�b����lI,��f�0"������� %P.@�9B�,+�
ʿ�O�䘎K�������k�C�L��` g�;��0�����r�˂gJ5US#
#���C�ӿ��׃J\e1�\a��op✉`��ʩO�y��~�
Y�K��B�#����t�S%Y��$���x'P�uW��mk���E�x^��p�9Y?d����ɚ� T�B��ZN�)�b{Y�[�{����e�d�a� 019�OLg�C֗���آ³M>%]�xə�v�Ǳ�1�B�r;��=�M���6�Ҫ��?���;�x��&A�Y]�-�5��o��l��S�_��e}@���g�$��)��M��E& ��NjU6�~���(�>uA(�w���cdR��Ur�� �\���i|�<v�ߺOE��Pw���6���Z̵�}�ނ��>��L���*������f�����or�59�Ǫlwe2MF��0�;��_���	�h�A�/S�%XqF^�m�N�.N��Q��S�")9�4�� Mm܎R�u�G�3)]��w�jz��~���oi*V�<4	�/w
���f����y��.�:jyV��P���ؑ�C
rV�N$br,U���aN�2�:d!�-��_}o���#�M���?�/�X��sCO;�,`��K������D�*_���w�rEvF.=�Ķ�;j��K����P.蓇(	;.�3�(0���]���٨�C��/sK�o���;�k��?(�B���mFػ*����^n������3�?	��x8Y�G�U=�-O��'b����`̪�W[\ bR3���30��ȳ'*��X�ʇ�!I�����ȗe�t�M��'*�_�m�|Mʮ;n��[����T���
�(�>.(�����0�J�E�Eua�Fl@�k&�(�Ҋ��.��d7���w� �$�;��&��v�N=ҿP�H� nA�p1�q�M�ZY�=�������o�T��:�����/�&
�F۲�&�ii������Z�Q��T�k[!;7qq�캢�J"�$����&c��2pH/�����������>���"��S�B�)0p$��\��q���@z����L\]	ca���C����}[Ym�tx�
�����F:��C4�*�Z����x�~������7aU��a��>r���o�>Ikl豸@ey�L�F��g �0�wz�6�C�˧�0�ȃ�����?O���E3oq\.�7���q�}$��ڒ�����TKG�OEyJ�����а����UFnHUa��}{x-�)���z�i?����j�z��գg���F0L�y�2��[�Еw�BkW&�?6�u��g�,�����QN��G�~�#�oR��:��ݜ�`�Qg��)z��
�TB	!j�/�5�F)-̱|4�Y�� eu�H_9Y��|�lm�B�g���_���H���?�!�m�=�e��(X�1�t���:�kT!�۾-z8bǮ�����Ab�F3����[pFP!��a¼-�	�x��F�O�p���
d�^�Sq-�\r5���9����!^g^hnf��Q����oXͻ3m6;�D:z���զ�V��+s�3u���\A�w�����xQ��<ˆC,��%D<�u���$�_�|6�MB��L5S�(Wl�]���
�-�?5�0������4�d���DG8 . "|Ghi�q6���]@�[�M��?N<I���� �gm�P�=�\�l��G"�T�q��a2�I��{���z�-m���������]��D߬����B���h�a��Im�+hU�3��&v�H�Ax��R�l�Қ���g��7x�G�x�����L�,;��H?o��9M�0�Z ��ݾxU�S�	=c�d '���.0S�4'�@?��֋{p�f�N�lV~Cޗ���c���Ǘ7Cw���(R,�حb6��<fӧƖ���j�)~�-�	�.��Ӹ�}��Ck.و ~����N0h��d��X̣�c�CE�嚀�Q���4��g���ّ�Vfg��/�|���/
F�g��*�L���Ʒ����>6��i#�s����<�{���`	��a�XאGU�=�^r��x�⫲�by���2[6������[v�j�:�O�"�¡s�k$x��́�_��z�� (���i�cL/�4���o9����^8�LF��X
�&��%��@@P;<�_	.�@�!ޝA�D��`~�Z��)j8+�؎a��fԱϥ�L9���`��}&����p�{�+*�4��kx�GQ�U���5lN��JlZP�c裼3��1�� ��T¡5��.�ӗ����Y#�S�ǶFj[����%=���B�n��k�+k�l�;2z�?�C R�v�c��F;9�*��F}%���|qNx��R�񔒟0���>bF���w5d���	��E8�)�
i̫���P������F�E�2�:񫟕�4�I�_F'���YǮ��lF�����ƱR;�bu4h�ʍf7>�唣����㞉���_2c����_��0ӛ�Z)ò�d⦾�" �����^d��ÀA�>���~Y��'�Y�P(أ8O�0k�5�h�/]��d��o 	5�w>�SM��F\[l�a�;�IN�2�7,��z�(��%����Ѓ��AE }a�$�(Q�#�!�*7)]5�_��xj�Й��C��pj�B�$N3��/�*�|<���%������N�ԑq��_���"�.��_��U����_�S�	�J��aME8T�(S�kb��6;c&?�u�>�^K��|W�ԝ4X�����E�VlA'�B��{�DdS.�`���Pj�6<��".3+[�A������Y�dzk��x��:�z����,۠r�x�o�����Rw\R�u���:P��Nγ�g� _���E��m\��t~�;7�ad/�5�����`� ��§���$8螗��6G���?�qʛ�m���·�����=�_rأ?��<��+�n p�8�t�a?Uu����E�BhB�H'<b�6�9p��r���qg�2��7���4C�T~]VNJ\a���=�������m �R�Vho�@9��H�m�W;��r����զ���TU�&�5cV;���n�� 
j߬(&�h�!��l]Aʣ�L�L9ofV	�L��u����F�aG߾[��=�'@��]���M6�h�Fa�d��W��`�-�ax����
�d�ԅ��ڔ�P���^�w��Z-�f���P��kz"����^�G�X4�hݳ7����
�g�s�W��.�իr��#�2>m�6����Q�tV��� ��I\�Ƃ��}�Jt����q��}��
5�V���1�b��E�:w��U5z=a�R�De����{oȕ��-d3Kws <)iޞ�����| �O� �[|�e���Z�I�s�����O�ț*�d��<�ۋL���o?�����֯��(�G�#:#����I�j��SU*Җiv��A�-e�jE[�a��mw��JJ9���{v���4��Z�]�F�\����C�Θ&�ܢ�qI��V�����>��~@h[kb��܅#*&�OWIL\g,B F��H�ͯ�5�"j�ch���~�~?��m���`�:E�S%���Hx���kٵ&���O����>����ӊ�X٘~k��^��9��x�O�/{k�Sv:YPa 0�4D������m2����
Dn�%Φ�:���2���8O0����\����z�������	^�9�S.<h8��[`=h��O��W��_=�jo���,i���_��F"\`ֆ��bY��+pUMrw*̃C���lH}�}�T2u���A��v�V�*��B��_��1��Eơ��H_LC .�٧�M��)��L���~k�Y7�R��|-��	xCtcR�'`��n���bI�;gF��~,��?9�P=]LEw=u��o��'� �KG��c*�e��2=1�r�q�7j2uEՁ ���r�����?vs�?C�ޔ�EE�Ob(�8v��j���e� ���ՇzLE�1<�b�M�n�,2�J��%�IS{��8�I����,�儡�r�����i(���}rH�6��lUs���OQ�S-�Js��Y/'���*ڪ�m'�5
1p�$����"<|�m��	�
#�F�nw��^���麺2���};�t���qS�+�U����I����[UY3dօI�=K�ihA���8�m�5q&��A���L��3��l�����X�l"���b4F�僝�w}��Ǳ�tE��AI|ƿ ���a�H�=�&yį �/X�@E����x,��ʝi��x�w�!�3#����TzH]C2G�Cu���d�fq��0v�����08C���iqq��T:��� ��$'��/բ�4�q�X��@��N5�]&d2����=��mY�K@i�m�@�>JJ׊�X�_����4���נ���ۦ��{[%�WPm���n�:fW*�T����:�**Tө�B����v�v�� ߆r �F���r�dOEu� �=��4��0&���������7��l@�/CY�J�)�~`��x��x�M���k�m�yu%A��jdHa<ڑ����v;촍bA5H5 nD
�\GNDa{�����D�I�f�7����RN$2I�O�Z+�"$׃F�7i�,.�P�ڼ�"�fEr�f^"��9��2Sٸ��t�|%�B���(T�O-�yk֖�GK�!���p�,�\`�E.�I^��Go�O��1׍�m��MR��\�W S���TM�=i�1m���#��XO0>N�x
�'�夠Փ" �ѝ��?�0'd��8#�:`��p�5KlA�~��3����h˒	˗��l)Ȋܰ|�=��C�@����m�mo��仳d�G`�8�A{ k�K޾��,��RzG�ڏ���z�)���Q�;��8�QZ��=�z����Q��,K�c��v��K�j����ٱ銔���q�П�6�q�I�i����B`�Rqx������V�O�y�	��Z��LH֣���������H]�~�����JvX��V	��$%3�/:K�x�mJ}���������W�����%�"l�����.�v�,����VS�<�/�=�'�CB�u��N�N��?k�.6��s���4���,���K�wLIi[�8e��߽��x�`70���^/��l�����hT��r%���D���+ji�Ԩxө��LA:۽i}%k�����^	��f�����a����}q�f���5̰���7�j2b�)q��q;��ֿ�A������X��8��W��*Y]1(#�[�g��"�چ~؜��""��K��ˇuQ@�\�Y��<��diD�BK���w1�7FTrv��]9b�7�E� ��f�<��OxEH'��q����OG[�͛o�sy~��8������4�ᗈt ;VݞF����&����8ܳR�S[(�Q�狚�>�:�+�ie
��:Z��ԧ7�1���w���&����D>�	7�uR�g:'�����!�;&��c&�$�9II�,ΐ~X�p��R���eLɜV/PlMGz�Y������4]I-�����tG�A�rg�Ů����~ya��;���7�y��3���͠R4�؇���G:�C��x)�>��D��(e���\u��T�-mŭ>�2v��b��~7]Em6�� (P�wcN�K�އ%�E��������yPz_�=t��/��;�2X����BF���!�v�3�2�Y����������<(uC���N�/oXF �ŨA���x�� ܫ�0��
��qъ��:�7X%9����IR[9�!����|Ж�����x�w��0&���s��D_!�����jJ����N��➃�qE��"zO��iA�u/�1�����Pmk��!I�g�����s�I]���H�a��VѮif���v0��a������k����T5HG���W�9t�a�S�)�6��}��D�V �iX��	G$�;�r���bI��<<�B_E����Ԟ�ۮ��NX`y�5��1\���a,�1�"�خKt⩱d�JA�J@���=Y�\�~�Jx�j����A�S@ ����(?�#�Qݒ2�M�bI����M����O�bz�|f$��+m����h�6��s�m�jd7�J���bĚ��%��M��7y[��>ԑ�#݅��sB��]d�X5��ݨ���H��k��""�ް��2�3a��<��&�|r���2�O�H�>L&�@��ȼ�#�yA�����3%��)��y7��y���4	�Xmp��Ka�^�q��%�Ko@���'���%ؔ��0�RW�7�*�a��rI�'&��-<?R�q�}���{v�j�&93�����Z�G?�k��'ۜbU���ڝ@�X@C+=�NS\F�D&�,�|2�}2R��[p��,�]�+�XҞX���n��10��1H�k"���f%�#�]�� �R��hNCr�svl|��	���n���b�4����'�pF����J�	3*���X�����;;d���Kx�;ip���%�U��2c$s�U�00�{�� ����J�s�(��E�˥��_vJ���|@���}tXKx'�W�\��I:q���B+�zdxaa.�F`��Y8�N�[���Gn���M�;��K�G��-S�~���KXS!PJ�b�&�"|v�6#LŁ����ql�5H����n�e��=E=��'����F������S�f�mhRn�E"N��],������4�uU�@�t��7���;���&C5��G��w�M��/~sty+����k�[V�b���S�a�,�3c�F�@���Lق)�U���B�q�G�1����m�w��2�M��p��`~��g*y��Bf&N��4���el���u��Bd�+����`��Vs'�I��p������6^��)���g�_v��׉�'��$=�+\��e�����-�`!0Z����F���!��>C��o+_�?9�<{8�'����!�`�����@kĢ�f*�l('������z��Ƣ
����1�I@F����X�	R��<�'�d`�|UP��/'�c��Z�]# $4���Vٿ��d��X���8s3̉sƫ�� \�[:������24�?�1�����rXo�Z��`�4�'ؤ� S�&�s����0pe��0���.��Ӵ��wg�E�ҐfIko�_��À2h>@�L����4��3u=Ie�����?��}20g�%��C��<͛I^��ىqV��~eX����z�%�lpE!%&~�7<8�["N������$O���������cwE���AS- w]��r���v�H"f�:�gw�����3�"�A��	�0bP�"k��5v��O[K��ʋ`(�I�ͽ�\���n�UF�v2F�#��,��W����h��Q%���f�&��B��V|I︷�����1"N��Q�,X4��
�DC�&	�Ԟ5��˧C��t��Ơ(E%q?�)[�N�̫XP!4�\/������%'��V<�qh��D�,Ǫ�߸WXJ-_h�G<��[�~��j�=��eׁ�0Y�"q�c��&rEA��U��.1<�fk L䅷ȃ#�R%ҬK��d�xE\=1
�+�c�uMB�>�f�mI��g�.d���>-���8���,QŁP�>����.e�?q1���j�5��s�i�X]=�*�C�"��L�^��ƫ���v���*�h�u���2�� �Q��%l �R��30���<V_x�h?�(��;[W��d�;q�q��b����J���sjL�{�*k܄t� @lo�����ȏ��o�߼d�+��P���P�����z���N�?���O���h��n8�ǝ�~lG��c��8���q]�g$ <7]����*�kB���^І}��bn$�s�0�uҥǎB"�35.ȗdJ�>�޶�꺨�{wp�����P�J�4���(���c����J���DHT��]D�ҭ���D�1Xt[�f��(���)��OYh,��*�R���k�������a�j�����9?vկ����8��<.ey졷 ��(�s���x���0��'j���v��~I�R���SK��90O<W���'��̄��7�L���v Iu&V�֡�8X�JJ�wS��zӘ���)��S�e�k־����h��i�	T��� h4
�*��d��l]W���절�9��=�!B�tWx�!o���Hܑ�7�\$*����"�����Eۀ�G��f�������W�ׄ��9�I��"EgT�Ѽ.�ƴ� ���%FUCR;��Ƭ�ryk⾑iY�_�(�n�v�[f�>�Y�Ee�w�)ـ��ȱ툃��ZK��RsX��������%*0(��b��\dm<!lJT-�	1���mצr��������LhC���U�����Wth����3�<(�?���v��E�9�
'+���v����Eqz��s�j�� �G����4|���*���,�����;sPlf}k������һ���)K�O��+�(�{,v]0��Rm��f�mmT���<#.���[^��^�N�N0)�='��������n��������;��q��E7��l�[	Uظ�,�h�g�N;�11���WXFRe'�� �p�X��rf����Fhq���v�����JP�W41 Ы��|/Hp����>��YC�H�ȧ�[�k�Ǿ�u��������&8��͠*�k�e���_{�u
sI�o:.���q�Q�-WUZР�m�5
�N�VXd��6"�W8ʜj��D}���U�P5�:�:�ۥ?11=s�^�ƛ� i�u�[P��h��v��%���<���>�rzE�,��I�b`$í2�PO������}��k�XB.R�u����؏6�0��7'�s����R�����f ���ֆg?��#�Ň�׀��"¶HYd��MU=���wVJ$�x�w�o�?@�2�>H��G}��Ԫ{�s
z�~X�>��h]�M��tuZ��(�4�Ҝk-��*�Zx(�*W_|�m�U�v��H#E��n$a������w�R�D�k �Gߞ�:��ްO��^U��E㫳�D�X�[%{7V��#Ө�~����"]�tSd"h��b ���O��|�4�$64F�����fF�x�����t[�ʩ�r<�!�d]�H,����-��>�]� ��u��l�ѽv�f�8�_9�M�Z0��.!���E�X�D���N|�O!i��쵙��A�99u#tb0�OR���e^;���)&�f��;�FK��u�9�7�w����3_�9��ۀ�s���g�o�&��/r����[^�uo%��Wj��Gl+%�Dʴ읧��^[���EG������UL���#���0Z�9!�N��}GS����Wa�%�ϝ��5h�"NT�k��.Մ�,խ��:��_};�;J�z�MM��k��X��[�����*p֪;J�E,˭N5X^�7 `i��.�� RɊ��Y�eks��՟������|�S��#��zώ����Iyۿ��V�p�A�\� �C \�͈�pܒ���kdRTo|���8��x=�%#cq���[!�!�*a����A�6%����qs��HE����S�MQ0[P4l��R��I�|�=:$#c����[k
3���yK��ʯ���!�y�<ג@z����Lp�:P��5
A��+��V�2U��*�N�1V�W�