-- (C) 2001-2016 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
wlorcmTqaukoTnomNesgavceOGG/6h6PLCEujRx8idCfnIpZsXEsHhDmQGS5nyTFx4xGBgq7h/Oq
9KtFFYZONU02VHdnj93Bbiqea4Nv9wEgGJvoKSfv25SfJq6X/lvz+dB/Aa9CsCTLLWX0gAJrJpTk
96/6/r3Fi0bfvk5+5iw2NP7Cl0lm57hzabFJDehZI2b2g4n+jHdcsrtC8zbToiGC8RuCmdMwSago
Ajz3UQcq4C5oqe5crPmT3VqCOUt0oaNrE+iopo3obhnjSodf7rUYl+Uw6u3Ft1D/HXS+AcpiKizB
0+k2vVk1F/kAC+b7Zc4948Re/3M1uLNvWSo3TA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 16400)
`protect data_block
3PpEw+uMY1vQWJzkjAysRobsYDtD7L8hvrDECBEN4DG0/zDj5Jcxs+G6JKll4JtxGEqGNb5/0smI
GVhkinpjkIchYFunZNdPmG2zyounhIjT5vHkWPNJfAj4gvL/KQp6EV1hgOfRX5h8tGG9k3/qqGBl
TIICleS2f1A7bQA06Sc8uGdWb16wUcW5uHI9kp+puxodP8Cptkkg5CjXbjT7MoablbyYQTy2STVR
9egasczFClNMZBk9HN59FowWO+biAVO7qzZklD7bY84t/n8uTY3hErDhsnXkDzrv9kWh0ERi5bKI
fuIuniJ1Vy/NPe5VKIVcRKAoJyQ2CfrEX8NtX+QVeJ6L3Hwc88BM1NOikpEKXn498RW/Ug7a/U3u
m9KFd1JQh2TA0n6GRf+9zyRyzKET8g6kuOEKMvJ9r6HlkP23UQLNAhA8PfXqxfM5VrYOwnsXJBA0
fy2UNgyDIk5v6zoK/A1hipiGHvpW/0Yeu3qQAEku3eRND5Lbn2FrExn2HmCC/TOdV8QLoSKZ640Y
F6qhAbD1H41JV+aGHkYtQF7wNS4IlCqqODSQoZ9EtQbWvXin67qg1aG2iPSVvbPUJGzERDybMVSy
L3C+AXpwVZYkvjixvl/dBg7OnFGA04SP7djKskXKrVwj6lbqfWbs3hPwXc1LVSekhOPrB2k+e++N
iKQxweDWxbEs+DKs27axW/iHRz7VxjW4FRl7bBl7YULyQt6lhvia+M3J88dKhhTBsAQLylS3cXqz
z0Tz96BIz49F+22/bD9ZWvhuErQfBwhg0Nu+htgiqwpWbfLJxWuZjJ5vwPLMdaQIJxhJMAGl/Ci2
5dQmWJFkIWFatmXT/vT6l583azZ34QtzKJ9Qn5PEUu44M+Zpc8CZllKcu3m3sDv3wbYDYfnQEP81
xyRq04a832Q/vWQwb//LavM3p/RQe3g0QXu15ma1ERFiQKW+uLjQPG0s1feDqYHgE5DyQqCmo2qm
ixIYWDud7L1bAKZvuWE2/tVQJiUgU1fzu3I12u/SExulFJ3pg1CMbLOyYRe8yAJpJoRmjzRr/YXc
1Ii/hGwGXziDCvkpFFiDdeTVxta8q/cPunsWJDk0XximU71+Kr2S+8AlV6WFSQ+v0FycRltZQrRq
I9aU5C4EAM7jKONNbInwfDbIaYzQrER3If7s5j+zH+l8v6ufyHogNNs3+Se8CgS+0R7tQjXnMjy6
sO+QbRjUBrfHXyRppA5+J/SBghg1Gt04PF49WzQG1Qk0b+e2nGiT9Gv8ZBans005CDgov5KEWu5J
y18lg050jh5s+5kg7fExJ0u9246ttEtMKS/P26NDEPr/74QfnUUOXgqmTKWgiuGLzcYtxyaJ/x4T
9TQ91EvS6sbxoKwcBnjbPbZAwLZw1K4T+6zJM4rgiinnQeemyLXn5aE8JMNcTN8vQtjx0Oz/umIk
PWAf093QNpy4UHLlxa4kS3KaVzYAanmMEs0GxUzu5xyJIBDo5kRMU6yEGWTTE9Xp658G9I0MOLF/
Y031KkFjqv8P7JOBjHdVsRdBhfD/uYkAwHqFoObF6KV0o4o++df3A7OHYPcOPKywrVgePiQTVFFi
idJTbykwaOOQ8I5nVNxtuUH3A2t/aA0VDpwvDkO7tX9gQ3XYtE/tA444lZCfLUm+okSyvGaVnThU
Z7Aa1XVOvSWABTH5gwZjYs5AXi5dHdx9o83F9b9cD5xJPt1yiyNS71QNTn6mUI4SefDdvdmZoehp
Y16zca57SNZuV361QBuJME7RSHjuIj0QNgLXk45vI4GG2rnFCfYX5gKdXZiTfV+c1uxfGy2DMzAe
/IA0wHTdQ5luxO3ztXBTUibfeKlAe4QvwCE3rbImL3BbT2Qos+9mEszBnP5PS+cX/wrTaBRmzWJV
XQt7/QeYltSlStbReVR78/ag4Af1Y/nE43vCFy8zB/nZUgaW1XuLy2En/KzINCkwu0fu0WN4sNtz
WQTzcZQ/C6TR6UHuOo8x2qrfuO91RAxd3jUqAxnfiXCxTh2/oZeAEOJHTNwYveMyk/xjh22Dtywe
aXiWv+M9HlwNoe4KM5XPVWrGN/3yZHmzLLtHwNIs7AH1YCp/sFKwHDofkYrsbsOJ02V+XdgVvVkr
rqdiGnG+SwMtsWLvUqt6dBCWk6o4KIYm9PlFTKsF/4AE537bIBGp/yaS/76kbBn9N4i0VZZVuEq/
gkdovTEaEHTBlHVUxPM4Vtem+bF/gF0BZ92dRi8cBEPD5pzgHYcxznxXY35ZZiOGfVl7r9zy3eWL
Pv0DgvfAinW2+N9wPJ3te7G6ZNr1xxS8eY8zKRfCZ9+jNs9mvnJrl7bzL4zfFwt6OCvEwaq8b9Xj
W+ksBb6EtCd81LV1iPZFKx2PVghrxWDe7e0G1IDjcO0uRS6fHkRRsmyIoXTpdYRNDQZblWPu+PXy
FlfqImy02hCpyq6i2ymnV436kCGoyJxQxgo/7MQKl7dYbO/pPy/INJkVBwOVp4IP//MP4/hMYY09
vRp0dqPJfaEKXy6Qn+8XKz5gPlXEqHbGlSnTqMIvGYCjgRkRhNxkwfyM2QBSObpOoGJ/7+xtIF2p
7mmsyITOxzeBjtXEslmFfV/Tb9IQp1xk13fdKRIP8IKIIDm4IuzKog6uILqjnvnG0rD8spP9I1bN
JkEWahiKAw00wOhOXzhJRy4dg53EZA1nnW7tjQHDwtgo0rOFJ2/EWgJ/c1s/MwreMb9zLloY/8h4
OqmcTlq4T5xj7S4iLTNhkR2uNxCrTErE+nZJjrd1MZQAMrWQZgw5XXuwXvsKKDG3i/lQ4rc3MOqL
FuQrCMiKDJCfzBg15ZeIe1MM3mSyUTemvu+7Ki8CJVDPGPrVW/kwGf/8QmjOfo30NlUdTSpZSmHI
iS6R6hihRRSSOPpgM5pj2mj529IV4JTlktwD4XlY/Cr0NkczcHf9+vo7KTfdrDvW3flsU8z9XUlw
KoqzolzC/O4mLWl9olUBHbs+PVhwZ/z5WL44NmX8lZl9TSupWesm3JtnkLSAz5rqcOee3Vg2KsOR
xGXOtifR/X//1bQGW2nkJOiWOynaZsiczMiG59NuISvldlTzQEfDji0hpsOqQg2zAfz/dOH1BM3M
WJDi9VC5AxdNwo1SU3RZZX+sOM0nxADlvJ9I/F6QlnOaXctvg36of62VEdP241dZXnVacdIq6Q0h
mhATcDUjfJXCSqHDpMtL6FrUhDR1z4RDiF+PaXnkKzu8SU9/WOAuj8y3BRCF+QzYq0f4gcCtxEVH
gKpGu4DAHrkNmu/HD29aootML6lQHvNEaUk+FAIQOuRMcLNk9LUJrtJVC09IwzJHyNBf4VYYH/Hn
qKyESR1DCZGaVjjfsAd2Sec62QGzCK+nYn2Q+1aqbk+hCtYE1KhQptylcSK5MqAw3763H29TgGXs
K1atxYERCNRNdANncthjAWkUpeJX/abvbM1bIPRdhLv+k+dz7ipN1pZ95gyn6y1m8Uva0DuIkIva
mKHmwQ8cINkpQHPJLpIfnRPMmUqy+GY6lK3DWeroC+ntH4wcpKJMv4ts57Sdgi5+7FbAhAwojzgQ
kpcAoygKBe0RmL6ldDACZQ3RKd9WQ4VJ3ZhuTDAxB7SvqSjAnlx7doNUnIMxVSIQ+OlnX85KFuOO
oLMr+Sant2FQ0KykGCsDtEZmJ8tQn4uePnT8hYzweN05vTykFnjKjdE3YiZfPzdChLdpyX3oAcYt
mzSGRCnGDCeaTqHLYxNI5prNL7gqCNkgyc/FkTpJFhYEUC9s7FffdHgK0I+1VXYKc/GV9Bzh5qzJ
XLUmZoMdBl7SQe70GkOXqaCVseDFNAAJHjYY5TGTl3xqcVZt3XyeCqM01Pj4NPCZLyRhNJZzHAWX
mG7S/irYnYt3eoazxgVWjz7uoyEx4sV0jx5XX3GRMhLa+UazXMadpLstjt6y7ATCkFa9LgY4dcVL
P14Euu16hizhinKm/2YMMWuZplTvxKM3UL2feqAdWCSnPHpXRmrQ/v01FJJEhfCCwYDDRulxIJu7
Z/krJyBB8S762wFeHLNwQuoOhvD8Mj+IXudq/Auh6pY6DAYMdJl50jOXiJgD1FCbPzYX1BnsT/4I
7sDV598QCSSic0EwXWWP+RPUBpGgSQe5+Twnud4Yqpw7LEtN0yTvEaMj1GJuEGk+PXhTvogCxAhK
GPJhSsmpa6r2AcQa1yildtv9MhyekLREG3EzdrhR11x/VB/ld+/OWVazpdK8D4BSXobf+L+BNFIP
U2MlLdVxRFFXWkEri95CnlSW4CjlEHMYMrD1YWejbBaWdYS5Tz9q+Sa2y4YvKayrenMcQmTsm1ja
hTshCM6ApcqztSRAgp3Tfcdo9EiZ2DpCpW4aqxZBUaIETxpRl6xDnvma8WU8BqDnMne5YUNHPqpf
X0jk5/RO47sJzNLL2HSM+yYE7unNq+5QI70f5u6Pxynt6soAEav4Q2NlEv8rwxk9miRm3z4/vjHM
up6IwvJm7nypSblK53hUvPTlSnrjwW08Z4biVZYymPqIqgvicHiBnffmNRXEObHK7TYWHzEmCJMw
KLQNgdcLoOS1sksP5PKLWsBuT4sGijjiOUCNWX+LJLhJeWJjYfni5chs5iVEifG2iYpKmiN7tKUs
+8AKjPf89/OerqAzw9DGjILumZaSDHioX32zm0OoQRCE1YODvlCSQ8eB+i/GOE8LhTO2d0y3lnJK
Z9b+ReYo91k9GfIHUg5+5J/Fi9jkUwylCw88xlwHJH/0s8oj8xVZ7erF3okUiIZy/JDCQjN/v+E8
TDvtuBShtTT6o5rx8dFW096bZjhvGF6T0nPrM4I3YhtqabWeXtT6wJEH74od+vq1swSvPCNwOr0s
kRnaZwGWs8MnTnyQ56/eB1zM4uli/297i0SzBQ+Hvuo8S/XXNif477uqU3OiOZrfSgUqiyqzA3WG
7Oc4qhQIL7WOZwtWQbQOuT1wIEug5KYcFeDWGhVrwV8/kOvaJazctI7poqss6B3k4KrAo1ZORbsr
3iHU0dJeNalW9Iq4Hzr/YDseWO4QPi//3CqAixwm8s1IR9ZRymiCE8r+ALBbG/QKFwnGbg4evld5
Mq1YAph69WYIOYyT2LsOAzKUbnVHwCDPk92NrcOp4TlNW8mEOetpeJ3/TDqsXgSbLvpjhXPr+Zbs
R1ZqFezGs3qffaX8hC3stHVs+wDfuRjp0iCY5QhB4MNX0K9U1DZbqe+b4QyLNLuce15cOw/MnCQX
DYD93LsGYkPvZvKlF22i5mL0mZKOHxUtJSToBTscG4RPGE8WRpGVbCxCY5T7AVdFiJdghGLO4u7Y
x1uEjhyREzH/nQHMwzZ6NqB1uK/9YgC2csya1aFvsqFl8X9rQXLS89SXce17i14GZswwqXgJwtzA
GA8qSB0vqOKIcgs8+u6WCEKiTIqLqha16hD5y9QWh5GlyvO3b/nUT6Ilp3JsKB0EqbpXvj7frd2W
jB+wdGPPKZCDTg61ESecIupXoNWtQFVDilzQ9/3wkT57AH84CshlqQPYL7WVw7VbUQPNMgHWOIat
w5jbuEsASrmN8NFO5yUBCrPervQzts6oGlTLgJQtgwL5RFSErqLexWkkssAaevG4ZpfLRWinVtcd
ogA5//IdjW2AgNuDBk883oOCvQteq+v1uvn3QXA88/AGuzQwtplKmcBhLShoQ5pW+t9+kA2nh+Li
rsjVPZ308ts3hX6ZJa9bIsp2sHgq6bXOdDFY2yHAvrYYNKIcA8wJA10oH0ucXgTFHVUe4Sl4npMl
fs91IOXb67OBqwUSqOJB1Ky8DCGwr6y3RNpyVKs32r1u/1gzeO3uCTqk2Qj398BATur2cqXjPeTT
7yfV3mVVYf8tg/Liv6acBn7LDXhXlOge1GJVApKigYwP0T5k3/QYD8u2qKf71yrUO0LdzIF9AtkK
6v373GfnSKgrBcDqG4Kw33erSTVQbWdNe1ULuU8n6DTctkTWZvXgyb0aysS6KGgmikBKtofqI/Eq
FJbDfDvT6xNQv6zvT9G6rA02PpYIWPU7SyG+ZAe10nfObx2HnHyE3RkK28HQeqvQxIo8UfVJvQMy
9Kzte61M+x37QrpFiDZRLy6f0PYG1adlBk2CUc9gcWGyFwzh+oDh2/DJnTBHpzd89lI0P3srUyaC
cJy0lDCy2ciSATzzwCXCLbWDrOuiC1k+VAbTUZPHCqX7K4pRs6lrRFdVuFOP4dnQ1ESN0JBpllAc
8WVupeaYKt4kgE4TQGgnzU8rgUvYSzv7dD1jNPyjcJKIZpk4L60ARwCMoycFTmArq5eF//iiQarQ
zCB87mTu/123OGUwOTzS+niWQKiBWivlAQANZ5KSYIePFJOZmHGCjMNuVG1XNLvbt3+MJwgY6F6Z
ahp8pfII5bORWONO1VE3AZ0awxNT41dB5/EQD+hBO7qvJ63RgxQNva67NxnE0NHGWfSAF953A4UT
pAqGjPyEZLccXsnxViZC181LN9kJOO1l2fps3stDaQIrAR6DxuCBCPn39VyQFK6xJp4D0rJ6N13o
theY2InL3UNJLL8HfO2IVR6Q3o6+vzaPbuehJ1g6KZZWe4PzJdEn8dk4HP3nQNfs9JvuWab/Y3TS
0UOYS1fZTyyY3vswRfJUbM1XANbVlm1SksheiifoQwFWCqsT4BhsAakoj4VZdeG7iluPcqH0DC3T
4rrKWkAquYvFyPKZR3VOc0oqwRJDAlP0MF4GmaFvOxDzV5qXpEYv26P2OsMYwm+5aYHc74ltXgq3
NDsjsB6rNv0Z0YMiQNb0qpH0HjrNCzRsCVgL18825xEMdot9TgyUutcFdxKcgbk16r0pP6TCjDJX
mkF/C5pgwTWGfywTRlY/QWeDhmSdtdiCjx3+SUZ4t9Ufbd+92+aFZ4JSKBmRPWAzpZCK7GFFDVLC
Gd63Zg6NUqT04IJ3aPaVgiVJ0YaPndR2/9DXNA1sXt5Gx15MV/a4ZZ7cFMmB0Hj3yNyfQUXN4onO
fjBZkdIR3vjXTYEsQUwrQT2pROJitGK9hDV0+Ec6UiTKs6wp6JEkZZfBljlfSSJqreUXrmkuAtI9
D4Amz8KtlXgDtTAFkf2NolhXzCcNRk6/ptydmc+Eol425fnz1BunNJWUTJ9Rd9HtSGz20tD3Ov1w
RitHWL9rf4DJhGeFtlc4d0lXLvXtPAlMQ/AwsNtsZ4dAYkc1ClNVHYYTAfnZEwATfDRVPfoehVnt
nyCDUKr+qlnTrgPsjuij08oINwnEFCYUCMwSpg57zbn4qyFA7o81V0mI7ktCHMWDZJbI3K4DcSHg
0oykRD7la/GQxpVdr6XVHvMYiLQWqUE8Dag/11lKmdNFCUoozt1c1Ehfwe6r2LsOQ1K6Jtofynbs
cF/ixAdrAZWn/EAbuOKSYTaR1iXQJpECBT9hZ0T14+JSHWxTs1sbD+MCNHO9IyHcLLYerL0wwJ51
hbEZoAl6JMo3rK0kYOhM4iEbep7aqzowiJLWEBL6K0jGwm2r4+sDTCg2YDjj4K+y5di+snvh05Sx
BZTRFHcAGmSGG3E4Ku9tWZKpSXtkq4MT+Z+aYG9aRjHQOGDUyETj/m4ee1ojeym66nDetahj4J7N
wC3It93ShoQozpBuyYLqhStqbwJ3R/t4tQcES8jHV5yioED839MpuEvKx040kSJOgTX+bncILfnJ
w7JsoCVfMQX2E0Hg7hcrjZOwE/SMS6i4Rv1b6q83kbBDh82oR9W+KWsyon6fJBuZXtE/YV3QJ02O
O6ascTAlxpc/hP+Ge3Iad9KWs/mO4Pjvy6kMMa5yvvmu8EI2fCFdLrXSsEja29kJ0OeM0GeHIe0w
nSRxwq51SJgNyFICEr0CTK//HBxKb0Vi+Of3mck6x+dnbackOxU/XZ7aKqlNjxfROFG44l8q1V+9
a3115li4SMRTacwjV6fnY1kaw69HCUg9hY2JgcDmbBxIUBGwQz5lQIt52jjD0hT7VtdRzRDClJQJ
iASxp8a6wzNC4HjT+l62dyHqM+S+ovNPFvrwBOcnzO0SmfzQUMruVYH0KTlqkt9Xbbz7Plfc2/qV
tgNkSKWPyCer+SrZ8xAtSPJlIL9bKrZVY9ef18MwyPAzGXfViA8IkpjyyKwwp4TZAUcVuwAtkuA2
uG5+lyh+hPoAFlVVDn02CrIuGUAOO4h158cxwDaPgw4U0J9NkP3EpVciur9OoAiw9vrUL0+judJv
872Biy9O57q940Q2fUL62Z4iwbrjJTVIBjEbwUa6i9pvSGbduKDDSBtPrpzbTtGhUZfahu0ULlon
GNTm334NkenXmU3CIo4MFkgTbehFNu+stR3bem21uipv5Q3fldXbfYzbrQ2w7V5L/OwuNLSvMX+X
EkABpPUf9jNZo64S7WF4yNwmJbFpQjObtB19jVwAZVzxdgheX2Om60E9srh51yWbEZgYCowfIUwB
gW2SWeRzvDadicrwO/ZIM4iAqIU6QtjUMoLHVqgC5R73/sdDtAHEClu5o7MuETjjXoYc70yQQCDI
HspqxTpZD3ogoBaU2Nzow2jYOWLQXkNmk0XK2w9AH7rE2QFg9itTY29xDeMjbp7HLmnwdrpYDclE
E6283E88e8Thac6xflozxMdVG6ewBAeFKl+7Bfx8pula1ju2ysyW4utBYl8MpzbthSCucUNPlhXE
Ux0oz8Q7AlRTv3wduRthR1PZ3gBGNzfkJyyTKwZHLD37Kty4gTRtQzEQDoz5lr0+KFemymBZCg3o
SCWQExvMtIzaD+jqRLH9iyR/WSOVsq1qxNXfZ1o7tymGuCyS3HM6nUiHEfBoRTBoUR2gn1hTzwT6
lGnBJy9/VjczIeekEO3FiKJPin6W1z6kZNDs6QgXNUXURUY8oZH46dqvuZtaG3w9iYRJDJhPzUlu
dzLNgFB1W5rsdUQZCRZhdXJybdGqWh7GFR9qUQFpMmVO3Ax1a4gx6qUqT84HSC79hvUPrd9+6H+T
EzX7O6aNWj4pbBTJxG26SMS8QVoCn33ndr9GQzwntJX+AdoJvNmKLiNUW1EHgVppY5U00GK8ErmW
FqzX8ldtLO/BHRzmSQ0y7QHrp1zNoiIuqL0iYjb0LL5RvFUkgDxjyo8JYG4cCUskLJcQFFxOGg4g
wJs1dX9tA67L/gzMHkQOOyD8rV/NSpgTccWEMbxR0ZJbtqvdDocNC2R+qe9MUcxL5ETtEsBqD+Ar
cIIGA638ldLsmXKNG6kqqBvKsqkGdST8RFlCZHtrMyuB4y0qbffx77UV06JFhl2e3waItk8ppf/z
GHfmiQfDTzOpV5m7rHdbozQqDIA1nf8hJAFLDrAXQbmbtNaq5E48a0HlrTnkab01edfmENFf4RNT
OGz1vSNyFzoF3wdL6A3JhdxjTKnYvXyonD+1FmXYPM2/AfKDQRRNlWzXR91E/6VQpAORbqqDx85r
PQlhjfEzJ6IANOcurBWDQDvRrZkL4CGyt6T0/Qfg8D1DXYhroJZJm01v/lk8ekbkMIrwR5PVyQIm
9mRFMmORVN68LYeWfH7Y5dL9/L+TSGqNFVCaqHfjkWjZdZ1osUhOYGlhKGL9GjbNWOoXKHCkGOJ/
eIQ58ftlMdP004GYgFutV8u8PxgUWnUHak0rl9ELROUd2REEC+C5YCF8zMzrgulRXw8ED36TBpHF
Td6BHWRva1Tsm15Qvk7+bjxJYllFbYb5+RMekz1x3OBIL4KODObaA582lPJf37igeAw7pKA2ecza
QLDggsfhE+O6d0AKnGKj7JKtwTgWFNXCO3nhJTAp1FGunhnJwAsm7RqexYOugIaJvSJhD2kI7wZr
MMpVs5nOdIGMrrBvtcK7fFE7x1bIni6sgW4n6+d/4knHCCxsMhvjRHVVcpQs8WHcWuFNVazO+HGo
gtuPSJPmhFtclJ5x4eyCY6ST24+7O4MjPVpOEEU1KyIoIEcAjKzexS6vq6l/zKQdHEy6HE5f656a
sek5g2vIOJgPh7E3Vxj809xC3fgrjkYTHn5kqNDxDpvXx7Qwjr2N/NtOk0U8d1Czw+/Iu9/nkXSi
y2ziibIMEVYDqwEHAerylVQ+nJwdi6Vb6PeJMvpmtMmMS49I4/rHEzB3wWLUBTsF+rdCsCb7KtaP
9gK/aqJGdrS+Z6Z9hqwDWxPy6XGOjolfzXZh38SfrER3YJLzFq6JS+dCLKQfDFSwtLNsUocY0+9t
WLbbGzDpZg+n5YQsPGwEHnPklpRMqhAEFJRY/YjlPGb0Xw3g67RDiME9ZW23fY5xa/4zYfblkzfK
8QuSBLpG5ATjsitN3v2QRx7sTxGv/YEQryMdrcd4oLD3CphwzTY6jR4eORi/E7Pharfob2WFI1/D
E0vkdAQfR4eV0H4WsVSV8z36arWhfpFnnXyytqDAXkhdiY2NpycpiJcvR2Nqol3YZnF8m5KQueuN
UvGTU18aJa755dZpg6DK2NbeoYLZmgLeO4nzphIYR6grkwDzbjSL0yUpj9Q93auR3jCpyU2/HLex
7OKZxqOXmBMdlLp8wOAZEhqYEbkS0p+TxGFaqsWi6iO0HEnjLPHZvrDmEJ51GuD8Y8ZEuGV56dX5
RN1sApNUDh3glKJfxnRpiV3bo5hQgY4F2KAmvK5fq098yiNzWhLkMuKFGcp4CvhcjLpeJzvPeR3F
R6BKI2FBgDFq4U4ZbuWUksoEiA9FkblMAZ5TyHfkFmjnE/u0zzqdwDA8BMRwKgJHIFyPvNkCnpTP
RF758BIjI0XbaXlgQLeR9zpRdGk5I4LSButMNdk2pE4eJE38GxfU4Ee7JKmyL9UOTR+mLc5yFje3
kZ+JNLvgzYbT0WnjmTL0XMROzVBqS4zzX0ggyT/9eTUqlrD30ziHTZNl1C1F06qcB2y5AADX769m
aAU8b7lX6RKS0TikdgEfaFh0f6744M2LDvAF3N35PuSLAxZmVAkitty69ZLeRiHqmEVG48IrT+ug
hoMDipgAgp0UbtiaEQMP7RjHg4woRV7mjXsu6pLgfJHuzRHQ30ySM7znf/HxFqApDLXNx5IGl5yD
jbEGQ3jeBXV6l8SikxupyhH+VR3zu9F5vM/XpIqmxN/OeTBLWykhbER7TFsrJBn7gqVgkHC+fvei
4TpZRq7iB8Yu2OB5wjnj45ClpjffLrHlMJGQ0JrTwifmf09TZzju/u8r2AZ/tOuZWkdZqFNZcuaj
HRPr3kBj3I7fW2Tez0bJ/Fo4MlMlJbd/rsNIgiPWoPIKqiNsIRxZGQbZFxu2pf2JseLuUxOXkxWx
RbnDoBPBXitK6f6UJuoppnkqearmHiR3YlbMc8Ba6vadOZje2ani+KQytDsOjMAtxkVt2WCGiepG
lxNJc4+aiFCu5KxUfwVVBb+YDfi7Vdl1HTIuyZvUbvMaeeHdpLL6PW8H7M4nfWPREpzJth4vQ9kg
5JiXPaauX4uSdnkqHVNiDinBG8/NWFiJYCURiqyz3prSLezAn/sgJ/UjV0BXUfOY+C9LVVGDNfZ4
M2NgZyzF1xJ6unQIerOkaS22/lzBgrXBKxjm8JzrjjI4H48FZuvuHb7Wf+yvvRG6FlBm760Aystt
ZJz6uCogHjtXgkEuOV49VUWyWHvXjDAhfmHOJ2ztrKBknm3mbGUup0MW168XiThDf+WSCpSodlpW
yBdgj383mkRYflODYDC9f20ntl4LxDvF+Dw+fqdzoeCUuMdmwLmfVnzoRQt31MRMO+QQKO1tdBTu
SIiLvByiUtElgubfNXoX9eeFimv2njfFc2lqgaQJ+/Wzs58sXd+OTmLc0AL2q5tPLf3kLnFdqodi
kyfH9DBjkVRazblJw0Y3RuHp+OjOmcsGRi06cGZSIRjFZYdfHrAIP6ZZU/+uc9Nk8dJdahkqjNnM
qc7nYgYgqdqsjNi13ksb5qt/iP1qTZs3aepK8zE4cJz8HtIccxir/9ExZdcCxYzjoId820WQkNgH
wMWIIt6V30psy2358rJqwMW4Ylb5R/2+K1T6tH8ktBuNE+TCl3QdOgfhtdoQJCpmBwKQTyKX+6KQ
C6TQyBXG3UmKzvIglEZrpMrnCX86MeI66ORHm7Gmea1eDMG8EmdVe2jMmMAuFPomN7gnKPbmupkf
K9yw6mijAtV8RNSClSkacWAsH1PyRyk3F1v3AzF6NjP0FMQwwKrNDbzOM6aovrIa4zlJjyrWcWFi
3L7qSwPReCLNk0E+giNO0sI5jbYvLZ/q+Tj0JrKY9/RC8QsMwRY05l5gltXCiYqQYNpE6BkRYS8S
AFFRQD1BiduVO6M+u+dQy6A0YakbQFLF+uqT690hVj3D2slkZOZEXSDeCmlNfGo5V64G5uQXotHw
GdaEUFtzU9tYzSlvTNI2sPwaRnP7jPdURIWdVb6Sjj6nh3Bw1IUtVjfj23uxjv8eRWqDP7vGY7G9
kcGJ5fJbRQefK7Bnt/Ug4ohSr90WWVQ/xALqbjrPXbI3xR73U1iE8QoTXnbHSu6VZERSjunl5F3x
i/9kzsYQDP1q5hFvQSVw7caXfxVpU5RLlg6TbqdQClX9DOSAhX6hZsaEBAZ/5A2RJeF3S9ji0Bgz
HascV90Z9ZogZOSG97fnIz4KBCdGBPqA9HLZ+M44lP/5N0WOqHkbLJEepyUKRjW3atl0LTINUaZ2
ZeCZUwDUReuM9h1S+t/BEBAubT1ZLiPmoZQAowFyp9pwiJT+4uGDh1RvHVtADYejGmJtEHdKq7gv
8TwHNjidA6ReU13L8fqwjcUMAL9E2VLzNhGaBHqF6t5xZisat+6DdxpNqo4FvC4vIKu+vX3dXVbK
SxoPrwA16+IrmoJyZri8QITaujtWqphcf9RCj7pFBk1gCDoVwHPhRmHhwbc/uXJIDqV1fhs6A9UJ
QgWMGc++QAw59BLPVNo/WBDUS6/ihIaNk7ijSA+XomL6+AzblpqzCz1k7/HI1TwGzlZRJ1T7fgft
aSzGA6E1o4O8Bi1xpGDbc0bpiLZTo1XDI0X/vvqZRxUgoME+xNMf7qwH0kg/evoQ606Jc0xwRl3p
LQeZFMHJPmVGVz5J26h1HAa+C+JTkM0xrBusiuvLuLuykWmkfSU5KVT5TUpQAEk4aV26BtUuELOL
GS4GZfPH8ORk1UTMmqEoSvvcZTUsh0dLlWSDDPdd65ildR+OSQXNcrQmlsWGHVoseQ2nrorPA/vE
b3d0xq3omZGVp9FchNXc8axlvOF/6b0+3Tw0AN8KMIf/bVcfouilXgMS3+Qoo8ICpSIV49pzkii9
LRgOLT7WY8d5j5Uwx/biWBhga6c+OSQ0UfjjAoV3jSaeiUQrgjkK1DIWp9JQRGdXCEucMkCuymLd
Ekr2zAtqjoPJ0mFoSbRdjSrAdqRwbUIo0nN2XJwGW6RXUb2NimpDfEt+KVgbX5cFQF39xWcaNDvg
fTXkL0yrITBrCfZPSG9RIjOrfU5iq0NYkhlqFU+VHWaOhyqzgqhmJ4S4H26cmPIRJuBbdi2gJfc1
5JCvP1F8yRZLQeWmEMga+aWw+4pq0M2xvhBGi18oDvlWUXJRId6L7KJpWf7n9Axd20wl2tmyrB93
ISoZPV4dSj4sDo4fxFyO4HEy29olZC2U4p5sEjFhW0LmEr2eaQ8OqQjIMXMommRQni7F1Ha2OohF
G8/JD4PA+TLdP2yfF1M1lYulU2Ol9/QH1jXyU6yPl1rtVTotbBWvoo6SElWBQZ1OftM7okmpp7Nl
aaOt12JgdIDXr6bboQ+PA5F1u74IJtsqoGIH4+ivmTsaa/FPNlVPAnq5VAF+lCYhwjg3H9KyByYI
kAQDLh32Ld7710nsCgnPdn08F4SQ4RrcXJUHVa/CuRJaK3eN4TKV6zb2vPuJvmgpSf2BgsRmLXY9
cSAEa5VQ5VuzrfkecFdzNNdjeXwkxD3ghORNBcqNvZPyaUe/B/eL0PzfJvqCtF9exwVUlY66Eh5e
Q90E4QuaTB1iG6U9vgZh2OODzqjErw9u9owsKZ2nBnLkX5KXat3cnDYMlw7uQcGhbXrBMMO+HQsx
QvfIXIrSW7DY370NHUn4svVaflrLFIkQtkBcfcLxLU9uPINajZmrPhZnVJ8FzaE1tBIrZ7ajIiNU
xInteEJUIORQV9RwJWNllD2rBmJVpqNWuwjpB7Y9klnsssg7nHbEdYhsmc8d/wFxDpT8YgzBggvA
ECeYUVhx36CwzBllNrBP1OpiKx98RAV/tgJNybBVnUKNbsfhn21CX7s6v3X4I/e0C3QFbvWqSQ6m
YsCmLtukcYsL+xLNbuUUMIvoVcsi4eySDRZbnRLptcVJrAf0da16H12KP2CtEwnh1QVOFV/Wl+6E
ARyQHOuF9uHPAFNFB+xJnlrBS6PxsO4fQzXOzLnnHjJ2gaiof4XnE+AxkU4KnGX+WEitXbmp0IPJ
ywAIBK/LOaGuufByiTvTAcGBMw8PuZpB0/y8LmTAqHG9L4NN1Q84/4y2ejPkmud2QMb3xohzPZww
mGn9r31zrsAwc0EonhkMHQxuSbu6HmDifanwOjdpTE1bxsSlHlMaUvuhSQGpkuqX18ySR82W0I7e
k7jRp6Fy06NcfLw/Gh1M/FrTETEDH53dY4UQOlYYgrzpX9W1dLON6HtgYlxvcae7GHiMU8gr1YGj
HIkRFMGsRmHDoxJUaUNm2+aOXmTaoLlOpOdMqEhfaO+SwWlk+g3FtmlCfI6ijg6Mma9aRIPJmuLl
3TfIqHdTbqKC53kUiniJ0FXpj9zpn5F8T5WHKmndFs++AtaJJXX9vJMYr5TSSgmYs0tyLieiQ8F3
0N0TAOY1BGSMv+6cCkVc2WKCY8Q+/rx83Nc18xmI4O26vyOISK6MokLZpVIbC0ePUsB2ENpysDHV
D1F1Dp/7SwsCuUD2KQVgDWFLMoDhzF+52ttYF37WLi3vuX+9pIoCED8+Jz5m/asVk8aFk3Bl2+NN
QuWo/HtjU/exXmvaSls4PbB0J/94k681NEG0jtwDGg2NeAJb6OViltvg5BflFdL7cTt7Et9aLs6L
YwTTkI5Qxh+96EvJOMFURcguBQoVYfg+hY2LKJvZ31lbPh0kRczXnQKfkENDAIrn7dNd7xHSBRLL
gBNIkAdbP0euxQylzBkO4PQ01ofMG+546jOTjJPoMd7Pf2U+v5B5AlcOlKxl0TEy51P/hcqn0104
Mbt1R1f/B2dC4TRZwPot70JFIB4SRVyzGdqEylDDEuRGHxU0CDVqz1ptEyB7RqEiGczLt7dVloYc
PsrbtJ4jloyhpaTKUMBLPoXwaot5MRlfbBhugRiZX9xa06tDgbJO6D3YpZPfa0cUn1gJRdmTApYq
v5eZ1LxkcabQ17KXrs7my6jownEsUye2U2zjpkj0QDa5gi8Ok2UG6bjYhdBkqx5PJIenJhB7dUIU
Fqidf+9E0rn5bbVPa2LifQNMbEmYDC1QnEsSaM2lEAQZY8IFTtmUjWLpRXL+OgOXEZIwvfEBtPhU
1Rvb2LvVPYTOarLaWe9qCYoe4Gt0OPngOex049phja9xhXJ73vY1OyffCRRNU3yIV5xYxdSVPVgW
nD4gLkPggaWgEOxmh9CMM7YZWP3R+JG/IV0jhsqyHrZs6Kn03fELG8451yD+ZdqpEz6lttEblzFs
5srUFg49nFtzKFlnCgJzihv1gp66G3r32EyO39xiZsDG7nrdpJOpAPhpZ8OddKgnzcYsBHxfkfPZ
g5GmusHa5WIGOjhU5QTRQdRODo5Dcps98c6RCFf/aaG8Zff7DVxAXaw3CrLhYYOisrUWnkKEPhjF
/xAwuYo5SPEKv2Kx5t4qxFVD6Qy/HOpIItGeJqU/N6T7be5MQ2nsVtvI0fVm06uxkvlV9+3uPcCJ
k+72U7r0hUTs9/h6SuDS+VnEHIiRdax6Ba2D4nMmE16u8poLzWyZ/xhR+VVnOKp4TxzjlMtMQ53v
OfSN0BLM0O9Q8N6Uy7zYI2LudQJSBtYrU2rUGb399/Xan+VCAxroq8kOG5p1Assnd+dsc8ZHyYUU
hsFb7F/IcjR1fvfp1qrvf2cNnXRrnGvwRpvb5S/MofOP3VmTUysgF+OfzhTHHPtKT+RRXleVYWpy
fXVrcrARyLwpeuZyeufimxUJdRyR68GTuh5HJqLhrSvi9vtmEoU2kGq8XYG54KwGbY1KmedPt33a
lO6AeNhLG3xIBnp/7DR6pUnjc/uF0+FhOI5BIjO3D0pcNVgwrurNGFjGpomlmDFQGlPMjhMcHPN1
t++PlT6ij4mZjXgLxlvAhjTON2ouy/qICOzwqKFVgxtkbyVbicjSdIoTZrSkLLx7PkP5tCa4cjqS
9R13huDVIO5pPpKS7XmXToTu7mbbPyFZwD7i4J+Yku+uJkIAVgEMHBirKOEO5dssm+uvLm0meByc
xPxxmuJENT3i2i0QDcY2Ry9wNIWSrTHi/7Ge2bIJ18Fa8VoDeVLsQ8bUZTN75pbzQaJbf1Usi1lQ
lVEOHnL7s24NWXcEhSzYJgwong9xhA8LDvwSbkCwv1fa7KiJ4tVUiBmB8QJSw+viKszUS4jOyO90
jB/PAPPoGQ2MkOCXKd0tvSEiAe228ysjF2fNRAPOog3pIiZ2JexWcSDqO44evV1bUFgOhL56hots
XP5boI8WsWDSCdKofxmAwSYUC7C8/MEXblo449cPjh37KVPn7p4TgAQw5nsWZ6+IHA6rZAUlHZVM
j224bm/tGK0vQ/rbTBXC7mNiGVsORnMRTBL7x6H9vqa9Ps1pFkPVZGZqQ8qHAL+UbZrVT8xXbtdb
+ldq9Upg6vWyrVXs+X5lWi77DAWwbiXsrgcnxt0RYWx4oZV4WN6uk1SmT6FAwrq+1/RbaH+6KMvL
xncnO7MYY2hrl+agKIy8Ggiu+6hU7q+IROE2Ipa1xhPunVMtStcz37ad7aD5j2zW+K+0gUXH7sv4
PnApfHQ+V+zKlQYrWir+SmbsYL1I3/wZ/o6IC/EMFKUkPKGms0ik0Mhv9KCkE8Kc3jEXHnagSABv
jU1MfU/Yi2ig0wzs5uHLyvJb7CNzrHI7Wu4AERmP7YM/qgynP0Cma9uEAgyJnbsVtXanXlAv8vSG
EDkEQ4VgPux5lukJ3ItDJQwY1pjB5mUewHZ5tfkhvKIs0vMkNCqY3nY7Y/+uF8yaGmyaVB1yXJNL
NtdX+Bp5SmcuA6hHuPcjEWPsBD5zlD/VlPblJHVTusSLkK7sAmAnS8rvyZh3u+qA8/RAbkf9FYTk
uoPlwbK+Ar1WF9AutZxKHaH4yZWFwH3gCH9KlmK8IPguEYtmAabt0Qu5wDO+CG7ICfpaQCGUfHfU
TlB/rfX8WFXOpGtELW/J7KJvYBEQIJ5SAe8iLS4Ikd3G0kr0K/LYd5YuHnoGVtQd1h3iI9L43VPH
b4FNvv1+FkKCjM/D2N2cNIzsXyPhfUJlagXW1hl1ijHkZFN1ljqiDAuoOvVqkrkx/qMM9JCXKQHi
3Du13vYNnpXmw5nf1Ozv9BkfJNu9bdU4B60nhnLXynoJ/kd4xG06bJl1b57SfapUdIe6F11ch8Q+
q2Xes//YGISlGzp8kZrwoPbR7hqPb9rlgs4GpzZzR6eLGQ6tYD5eiooVrEI1ZSEoalp22rob++EH
5Pcgr0uMG+ivPJkx4HCDztbgw0Tftxrzu7j06Jn8gH+XnWkictMz5NidoFtNNQ/E8ikbSj62ZjUN
ChMFNjflAuN8rQkYhOzl2RDqiYt2Gqq+oXxSLfpPXMd0iIXquzAHS7RaK/nTLbMGyosmETwBpywr
9JdC3vre5g2E1YAWB/uQ87I8iizJ9PZz9/hg8ipZ4rlglhxRezmn20aVlvQDiRlrG1ydhGomtM84
4tlHER85XE3ie7YELEDPxnT5Ia4PB3SOEoCxZ47kMOjmrbPRLAlHZliabaUetzU1FEr1F1UHO9XH
9coa9nbXTSNjcDfRO26/xB6XoBuMQs+yrkov1MOt4h3oXHgMFbzUofNGg+topK9hnAN1syTFrb0m
xthhiCCFmIBkfoLa6YoYpji43WZLupFiWYpcA/vsoyFBAhxMEgPyFPHlUlX9i5Ht5RJ1lL5PD4UU
9g70yIsig3EDzGkb4/XeZP5wLQhzyfvezPxrU16qaXOdWyd74yiANmP466gMxVHbK9uzHZiDy+01
zaFBP6nnl4x6L32Mt+7K0R7FqPnaenR0iwuMW0dZv0SHMbzRfCqOvqvquCAJk8qXkh6nn5WdOHaE
2Wg1u/Y/7w1mLYFZWtRY9GYnMmXod3ivy4O4T7c7ZRU874SfypSIN5pw8F9QgITAI1ljJrhrfJrt
Btk1V5luIjsWlXwSqjqY17ZX7P5wewsXeUMHF8YzzANZW0DN6zuiUCeIFUnGNfA6dVq0qwZ6ZW2j
TpKhJX8KfcWAN3URS9H8rVrKZjtusQr+QohZI4FgYrPUGvN/J8R71XUEeFAk/Yr1M8ZcylXFjN/R
eU3DwT1Vh6pQ36B2N/ShT11Lwigp/UUP4BIINs2NFHmeid5jiVPOU5nEvJKDV6V1xLxsc6/xUNW+
XbsN7nbe4oZtG5JxunSi2s0pXIFpLyzPja3SWiPBYJjCYqo3WKgLkPZI4Xyn+dwLpv7/ADyVrmlD
ewuLVtyKRP0jnsXqRVDsjBTSi9A3tixoAqicVBhydOoYbJ0RVmmrFHLAJ1wlWOm27OFeMiDED+PK
ky+//K/6jlOe/l5EZJQLHtze8vOwSTIvHo7Hu+V2QzV4ALI07WtRs/upzAf8n+m+F2olDtuOkQJr
SOMhdpHIQUgU38ND4TO9MG9J4PqYmJ07ZXhg0dvtS+c3K7i62TMyvJui02/8OIDBZVsl70Ezly81
iNTmfsUOSy+nOnaOF8ZoF/8tncvpgoeRKNzzina0d9BIK7JFN67i8kjLL+efuO1h3hSpXCb8/WUt
zim1G9EdnC6JTFn65bQIKgAFg1uK6bHWghSllTvOwVVPaV9Rej86yQxo/gsbNaiguCL/zUieolVz
IbdLiQFhv00X6SS8shozruqQadQ2y3XhAusvQPvzmcakgFrLHW+Ot1FseTDYEef1alqs5rfkXITe
I6Xs9kjyMdxWBN6hhlbQWnO2RV5dU1/Llg/mpxna9cS7hn13KmMJlip9SlFCpqyZWMcw1HDDKygd
qul5z3AGJiN3s7sB2OMquWT8bM4gfTad5dK0h3lYHq5IZbZA1lqvVa0GBfgJCnUybqTSo5gTr1wp
Ta3gB+S7sGCxV82ZpagTvuyrbss3uwWEuDypoLBLoso6Mph+g3RbKkFCOyJNL+6QRUE/97f0dNQf
6IoyuKmLhcdWudGaayUQgOWcApIyR/cZVtsY7BhiCDrElNSM0Gpny0f3bpQGI6hwzC9y51QdO5a8
jFEgDKb6vvdj21EJf2Fongcok29eA7kj/o7O2A+JYGQ2a8xRPi/QOIr51hmpNTZQ6/Z1HDBVZ0lq
Rtse/AB2J79nLcmYfMIuLAFyeVPAVcPLlGA6CIlBaXe6D93+tJpDcmeEMvJ7lF3hNAnSx56nnF1F
nel06przWHBtaLXlv43aHGZ1SYfm7P8Qgi3tiSATPw6SHYVQI+hqD7xmYC9bAFvHFO+XPB3OQXDH
jEeqdtyAFgXkN8C+aC44BnFxkfHp8M1LseaEwodnJg184xE4Uq/HyT8rqcR1PbHng20skrPIt19Z
m40vR5j/HK2YBVxrU0SeDtRCWK0v7+OsTGwuYrktdB5lGPJiABSvvFAyn3anZOgNbx85D0l+0puv
qFiNHLJ/sNNYPYaM1fetCOgHBbMXPuePVuQBuxPPmYQXTe0NyNOT6a5/y87905j5I+zHNSxZeafK
vfIO7LCjCLgiTd0gH3POuFfJUlPWXDkm7NZCY/BXonpOgoyih+3dd95W1UhbgU30wtnD+CjGZJra
u+EbNtLtEGs/ROXHzs4V7TtvLW5glBUsmw7lg7a8Lu4PpDLcGGeE1ptSqeFOdgH0+6yhOzOHfJO0
gdeFylQAMrHFBOD5cAn6eiP2fGMOe7efrRxjMQUYoklHLNhL8guRbaJyVS7/t6pmw+NkbciTtYW0
2nmPjgqTdq5nO4gB/QCzlYrb4q7nDSTq7iY6dVJU6za5quFtIMsSuL+rncz3VyzHx7s7tyNzg6b5
3/y1GwbnJYbQOWinUxUCJP5aBcwBVMm/QIpfvLczvZWxxSCGLmQXj+FdxXq9b6cyEWTRQU4psmNW
ops7YHYQNFrbBiTczTfhwI30WHrlhc2kSKhgfmuuzNnqs9xIgLPz8bD8DNA5q1/2YgzXQT+m0Bgm
XJUtENDxiJtkcMv4nQu65ct2f6FLZcRU4w9IquaLESSqwg+XUwr6gWfcvSuOfw7/rFwq/YOzTYrG
ClMGkUR9DTl/2ePW8BcwEvVu1GNeZ4qrcJniKUYRloSNiT3JiN8WkBiMD+ZbW0+E84set/EZKAIQ
nzNUDESP8Ka+BiS94QSN5OzyeoDG4/D9TlwX1dnHe2PXPAMTIUcvqKybqoob8DtBmWUN6TxTjV2b
Oo2rmYopx+oOzZ7GtO/YnBNIwgsShpvL7bUQ2JwMcq5oFu3WmFDLjlCpyIdyCK3n7yran2gt2vV9
uJ2RM0CQbELJEI2HCTZPJCsAbrg1RJWyMe1pM1ez8ou7n1EcZDlMNPpLvxee3gFf4rFabMlwXC+G
g5+WZY/QoQV/KkmMH6C7EG2s0rPPMG89uueocC4rdDXedRpRvQVWMuvIAyFtrNFNzSBHcGpuHKcK
JQtW4WPiyH+2wHUzOjKWmfhV8SsEdaTEpNkPypU2WR+QqlgE3lR5gTp267/2UVH7ploCWRJh2TG+
HDFd4uD25cWCNhCPXeX0c3MALt3i4tvUBPFw1X3EopTHhaOLqu07QuB7vgnu/046PjBXrZ2TQZ2G
MuIBqas3otTv7xlE2Tee9kwew8GGOSr9rbo6r3eiWHRV0FdroOEhu8WpSxRY5pkS0vBJYmNLu/I3
s54P1OSZ7c6NwjrinY+HsUAcFuX8gT8N9WxNuK998oNsdHtJpdPtoVa7pQTOlRMRO3C+Ry05linF
a4YRAimEnMDEf9EMuxXeqrbiR8FNDOfUzEHedrP5KTnM7fetYmKukhUdj5s//z7yYljqs9OUJOom
Xf2MkM9y/ovbnABbi7rhbnte+anT1TPiH+txXX12AzTeR5SMLsMDFooNZdICUwvRr34snzWq25IU
qWkJv0bEvu5Dzfg7apAp1Af/eqTZcDhKSXBynHgRpff8pDZuoBqTIrIR0OzVuylHStCQcuoXzlyQ
dvXdH0Zc9dEfAfcDJBuPuOKB5NnehwBN1Af83tkJAupoa6g2Xdu1LIAMuiM+MSraupbiaPkak/vO
FNAOEgF7v1xS55Kf+SGIjzyd+ERP6hULcAttNn3Kp4PdATkVJDiLSSENlmn9M8sWVfAKwpWVN3su
KhHUMe4C7D5aFbiVtbdkR6mJIkOg4cqtLsP3Y6PgfRH8741Bq98chOHZj/JDbLB8wEDwphGTWP+H
A5BJrJ7krDUDHYI94fQXhl0uk1BTn4pWq9+KI4OjgvIsNhVs5keQnRFXUM12sBBAzmEc09H2Xb5z
/U6LuO5n43P3ytK32gwu7ENTQgfPlxc9cbk1mPURGayWdlIK76E1wlcAEC/hmUBfZUM7Zj9QN+3U
NqBT9tVuFxWKz4UafXX2slOAWbGk+pI9PjxBxgQYOcZjEJYm9mqyd5Y45Dz4VbAkxM9SM3dkgSEX
XroD3i12YZAid+ZZIzrzihlLZV9YJYJehXzykYOBkqgE6y9TYHO/hVwZSbrNp/jzaSfs5uYZBv29
jBVXSMU/MZ0ASx7JAFWZA1QtpxQ0Rynbo89WHelUinsSIDx7jW1SAyt2bspT2EYBc5+T6hs2IgbK
wW599Id0Wa6g7v9iuhJYL2mavmj39AW8UnW1ZlIAalzW0wbktMU2A7o=
`protect end_protected
