��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��,�y�}�ǰ�=4d�H���`I"��W�`r���T:tB�T4D�m�)�	1��I�t��
��8(�8t>s)ו�."[�漆���]�~�]��;�O(1#5�-� 偙O��QZ��~rL'�x[�i,mׇp���O�I43��4d�,�H�����SN��d���3���r��m���̨T�I;uj2Y� Er�*p�Q$Gm���p�V�`�2^���,hz�<p��l�Bxt�5��s��\yq���#�@W���f:m��T�	,*�񞭋����_��㧋l�	�\�:��uGd��PǷ��N�I��_����Tuv� ���us�(H�~�{2H�:Zor�Q	#%�3ˠ!��iS��95�,?�.���/�F�i{#���Tp5����Ҥ0{%���2vpn���X�����@l����3dc�ק�3	�Ed&3�ZN O���z��s�yxӡt��v*}ԫy nj#��lc��m戭k[��5)�A#�����8�!�]�Z�s�M���t��w�!��'ÒE�rv��Ϝ�c@<U��\tq+��&|�&X1)C�����r�A~��B�&�����s�:n{p��͠R�X⺂L^��R����c���f��J^?��ܣR�O 1�rV���:��T�4���AD����˩�F�w��)Dm�O�b,�a���1$��c��7t[i2>�ޔ0,S���󧇳Ϟ�ᒨ�-��}�!6��Jyv�醊�^_�(�H�(y^����o#����X��3-�k\8�M�T�"`R�DF6ȕ� �,5�;Ҭ C�k���1\������k�t־9�}���� ���QHF��"��t�9 ?��{E_�7��!����](�S��0�q��w�9��=�i]�1�GʦȪc�W�XC�|�$��}q�6�\�\���Bp��~�1��<ΐ�%{�%�3e��)6��I�*�K�X��q����y�>��sR��u2��V>曛�aŃ����Ur`iB��O���b���	�g���<�%>�N	��6�K{�؂e��\N1�Qҧ���ě��Bk>����yPQ�Y �r�E�ϛn�0-~�ߟ3����7�ɞ��W�˅�e??\�q�WY @RE�Xw��J�� �R2e��% 訮�G�ڹ���ײ��D���Lա�^�p.��F7�g�ɳ�%���f�#* N������N�|�/����C$!���/LQ@�W�ol��B7Ae�P��2'c��S��g�C��<.��a�\����QK��׏q�k�<v�J1 ��H}�QO\���'�N�':_����^�iU�D;̖���c6{/��S�UB��	�z'��͵`�854�����[�v<�l�'��H�Gf���Z��I�Y�`?�=h�/i΄@�깴q������`�	��ެ �(��XY+����/`���D"}�^#��\Dyr�//��G�����H�}�."��6_���}x���8�R �[v$���.�mi�`+���`��2�]�c��r��$|�ڗu�
4$�l�N��ӏ��݀�����_M׋qf���S�v�`���u�+I)��������2Kv��CAH��E�]�s��_cae��]��<�)�w�����A��+X�?@��}�2�Z��	
9�!�{\\^S6����YRoe���(�`�Y<M�Ͼ��9("��(�s�9T�q��8B�j����j1y���8���?8��h�y<$:�.�:�;iPSsw�d��*(3�-�� &�2`�f��M��"*z}��ͅ��	"���M��]��K�jxet����<z<����U+$��Z�gb\?�H�5�3)��t��Ͽ�F�{�B~Gl$�.�bt�vF�7�J_��E�-��P=��s�=�l�^gU���T���j%�b�/��v��)Ӏ�	5ʺ�u�H�F����t��������bV7;�L(���u#�3�����4�v�����K:���g5������_ŒQ��y\���`�����ִrB=��~JZb,Z�G��$n���z^3 a�(�PX�Ǣ�(t �,59$e��ޫ�XV���x���ɭ��[.?X56:V��m���|A�Xv��	���*�Nmҙ�r�)�^�H��?�mPt�#���b�S=��$���_��X�3*,:[S�� �����	U�~܊J�^2k�*�qX����6� ����
%�^PV���h=?O����Ŕ3��8�.�$�6���GAe�2���$p��(����[��{�K@Qs���X{)p9��l�4c��tgl�����
a��h?��&в�/�N>��n��[#�V��V�n��bNf�s5_� qAs�X�zX��<�멽�n���4�r�E.-�W�� ��";���u����!C����7t�;SJ��
/dk]{3K���4��K����fGG�m͡���HՄl�k(�?�n�op�Ê[iNJ����(f��Kei.�����|���]�Z��;8�bH������S�=��" 2�:tH�� J� �xEnn�^�!���|n���ps.�X��2�2\��и��7����.���O���$ݳ���s��ېK���@,Ϩ��sU:|��	曮���'��άg�z�^S�NʰF��e*�ñ� �t�I�O��*�}�A��u��~�0��W���_-[�E�H3�8*%��n����dۓ$�y���A���R�+N;Р�a21�az���:[t���mΐ�豊.�_!���"�L��9��mP�ȷ]�yX�p��J��������a�Yx�Hͤ^�c%��M���x�a��F�#���<ڽ`�E�w��%��-��f]�'B #J�F��%�.�e�4:�����+ o!0 ᷖ��a�d�򛍚m��X���{�R#���{�N����1�n����AW�~&X[�_XE�ۼ� �h���� 6�O\=X	p�GZ��. �Ζ��������; �c�C6*��<c����)+t[$����\�6�&(/S�'��Ӥ�S��>Җ��)_���@��Fq��D8J}��F"<M�gK��
��%��Ar
�����Y`�T;r�h��w���#-��~͔v@�|%Y'Dq� �M��&�tIM�z-P:ͫ�%&��j�	�Ҥ�2�7%��~a��Mq��\r�����A�V��O@�/��>s�
*dN�rU(�� S)�޿33�Ru�4
?��u�K�[�?%������IM�t��Nvn����%9Z$�O=���	i�!�q&9Z�P1���G@��;K�ުrab��
B�%��4p�`َ�N�p���\�,�?�����>�D����<�<���uT�^fv��h��BSQ�\ԓ�{�����yH��_{�q�p�{0�>�1jb �0q[r2����,��5H���;��
��֡.�1��ڃݜ=#��[u��҅K�Bh[��ų�Y�EfP.�Q@x/+�r�	Tc�L��j,�FU*��ê��+����(�4���Q�w5�� ��0��B���:٠��jw��p#�X��� �3��j��\BeT1��H��'�7�Aqzy�Ę��:K��U*�g���~��8���2
��U�Z0v�I��R�=5�����S����.a�0R��7k��*������U/~*"���D�[��|�͟�7���� �A��M��najA#,����#�9�R��X��H��'B5�	�M���t ��������W2�Q��m^���G�w�[����Z ��x�#�k��r����S�}{w��h��d)�{![Z�I�9��l$D�$�c=�K��B� ʲ��V'J���)���Vö
����1䭂�TҥT�-I����j4GW�<�`�%��� 6����e4�oQ�

R� �8U�aS#,"E���\�"�	Uf��
�#d�2�2�}N�ԟ,�9��	ʨ�Q�R�����p����eB��"H0`r�l��\��%�c��H�/��c��с�އ��ZĊn܃*,^�����RҚ�7)+�����!��Ly���_��z�1*