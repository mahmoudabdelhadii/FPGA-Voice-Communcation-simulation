��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��,�y�}�ǰ�=4d�H���`I"��W�`r���T:tB�T4D�m�)�	1��I�t��
��8(�8t>s)ו�."[�漆���]�~�]��;�O(1#5�-� 偙O��QZ��~rL'�x[�i,mׇp���O�I43��4d�,�H�����SN��d���3���r��m���̨T�I;uj2Y� Er�*p�Q$Gm���p�V�`�2^���,hz�<p��l�Bxt�5��s��\yq���#�@W���f:m��T�	,*�񞭋����_��㧋l�	�\�:��uGd��PǷ��N�I��_����Tuv� ���us�(H�~�{2H�:Zor�Q	#%�3ˠ!��iS��95�,?�.���/�F�i{#���Tp5����Ҥ0{%���2vpn���X�����@l����3dc�ק�3	�Ed&3�ZN O���z��s�yxӡt��v*}ԫy nj#��lc��m戭k[��5)�A#�����8�!�]�Z�s�M���t��w�!��'ÒE�rv��Ϝ�c@<U��\tq+��&|�&X1)C�����r�A~��B�&�����s�:n{p��͠R�X⺂L^��R����c���f��J^?��ܣR�O 1�rV���:��T�4���AD����˩�F�w��)Dm�O�b,�a���1$��c��7t[i2>�ޔ0,S���󧇳Ϟ�ᒨ�-��}�!6��Jyv�醊�^_�(�H�(y^����o#����X��3-�k\8�M�T�"`R�DF6ȕ� �,5�;Ҭ C�k���1\������k�t־9�}���� ���QHF��"��t�9 ?��{E_�7��!����]���-�p^8�3 ��TLM��q�"��z�����`%F�zU��K�^�Y;FI�$�*,���!���w~D�A�]�#����u/��eס�yl:TJ�a�ȆJ?fgu��!0m�e�ӵ�:*���"GH!՝^�"VIk,P�;�L�L�aQ��$y6�O�v�y�&�X�/#��Ot��o���6��պ�wr��U.���8b�6T��y�=��p�бU�{�?d7q�2�R�v����ɪb����5��F�p�E�X�Ĺ�#dM8
��
�5�n,�o���R�:*K��03��HA�J|5��e&��U1���0D`�����>�x�l4����js0��8�I'^���������cϪ]o ��"�F�؄�&{���1b8\e�����y����<r��y��:�c���*�WGC�%B7v����g]�����g���٨s�U:-���lÇ.��ſu��Z�5����lbh".�=H��X�$7�����j�@���|��m5���*@�$����izĪ���7�Ș��d�K�uA]���ȧ�)+z������d�My[\r����{�~}�p�$�1��n���㒲kH�ћk�����ɽ���S��;8:>�+�39�+�[����o����E�b����݅�7�H�r�$ՔX�Fe��jq�S,P�W����7��n���:��s��׋��Ⱥ>�R����dev��a���I>�ze==��S�t��?N�s��7V�k�E��ܺC�_6wוٵ� |zY����p�2!\��FW��.��e�B� SJ�鶤�����w2V�� ������2���2� FaM���2x���}~�Pai5�W��C ko�Y��\Uڴ��&˷ݢ#��a�ԃ<!�o 6C��y�\Ij���sw�V���)Hlbr�F������R{�}�I��12;�,�j���ui���}\d��x֕^D���&�jN�Q�E�u���&�έ(�3;o`��������o��G��-��U�
	\�i��^7�Z��6{@PLLR���� ���`y���udW��p�FU�:C�>EjU��L��P��qfE�g�H���+>�3�8��d��]	�0�x�9z�	V;�<��;�K�P"潘�:N*8߻+BA5�z�V���@�X��Ѧe�T
F'�u@p�V�q'���zi0"4�J�.�Y�F��4k������5�Nv��؇-Ƚ�Ia� �<zM9�:~���/��bT,F��(�uxHc�G���(ZP�d�z�e�X�P�'R��l�1���M����P�I+�_3n���'}1���~7�ؼ���h��1���fũ	b����?�n��a��N鹅~�|f\m��:���'��h-�w^<u���K̔��_�0��&7 �/5:��yAAf92jڷ���[�iUa������<^���"���)#�枨���)-r��g�ޯHm2]2\8���}��|oW�o���ĚA��C��h4C�	����yBu��kT��΋�G|� L���w��7^}��#Œ}T��<g|�[{�XO`�;�,��Z<ՍD6A	�<�Ђa�7�ꛤ�{�:I4�@�7��P8Pk��.�k��6Ϛ;C�;m���:�AI�{������*����\�Hб�h̀Ob{t'?'$�SO��b�cΪ�(�{ZB�.g�慾����ܐ2���|_�!_���A����DB�}���!�k�R|��1�F}��ci����Ӵ��#��p����>����>I��U���)V���jL
s��Z�=�BZ˪�">R:1�y �:��,@�2�P��<��;��E��4�om��5�$@�	����15`
�&m'	�z&���|g�MM����^9��įtVP,��|��Mh�O�K#'b���3�P���w����� a�	�x4�d�?b�
mI��>F��k��*��U^��g9_�)[�R
����2�g3G�s��y	Uܴ0�u�XO��?Gz5n�Jo��j'J�k�
F����d����<)%��]}����1���2��� á�Vt��	͆������F�g�z%�F��}������)��N} ������LS���@��C��-��`Y`Ԗjߛ��*\���ޜsK;m ��|��c|��b�j�-� ��t���ϐ�s ���']���a����(���C�VBh�A&�L�����m`s|�n��f	k��A�ׄ�O�2b�A�l&�h�T�厗1M�27�Ǆ�������ퟴ孊~��+�7��>W�N���WmϩS���%#O�p=�'���+�:HY��po�~8��D5Iŭ���7=����X�cq��Ԫ�ٝ��0T�Kb��bbg���H��!k�Կ�Ө�.~^�{��{/�4�5��&��iC0$r�Rͪ�1��,򜹖2��*f��iiH!%	���l#�����%��._�U�w+���9�	�W͋�L?�'X���B1[��RQ�h�6�_P��X�ٷ��4�'u��ޑir�,��H:ې�p�%Y3t&?��n�暦y��
��7�L�r_�ʃQ���;���9�~�,{���|��3E
���r�4v������/�<h���n%J�:J�/���O�����6���0e9���?ʔ}5(���������_M�oj�ݠ���g���~�t�L��U$��F/y��Y��/��`oz�h�	KW�{\S$���i�;�e[���{�����w�N[�\�RB�C[���"Fk6pD�����D�M����:Ǉ��f�x	��Y�?p��[W�)��8�o�xó�i�:�cC*4V����;}���*���Z�S,�P�c�ә�2����/*� Hl;N�`w.W ��Gq��G &!|��e<���Wp�`K�k�
)��JK���F��:���	�ֱ�w����N�j��b�@��@`bޖ�{Q�GV��F��m�K���Ǘ_�5��fD:�ײ�M,�*v'?k�4R�1@�<�"�k�r���~s�xdm^Ȥ�2O�j(�nn*����=T �P�'��X�Ԧ����=V���:�h���`y�����	�]�E�iI��b�2j5<�	^����a楞��n���n:��c�mʵ�ŕ��QQ�d�j����
�Ӷ�[q�z��Ao#"��D�}�����[�Dl�T�k�c�()�jT+��ϱN.��r^���$}xYQ�4/K'X �0�Զ�<��=�f7�&)��~�-���{��⻋?�b��R�7��Epw�<{o�J#�Wy������������%��M�_R�/~����[����	�d��K��Ģ#b
����P��>��^js|̊%բ߷Gg�y�	C��8���rg��9�h�[�}I��M�s�b^���|r����8 �da߃E��Yh�Lt��������ص��'zv4&�Φv��ƾ䏤�M:g��J���K�K�>g�g������E&sAc>a�X<{)�+h�����@����d�+�})�Q�H���o���z�<���5���ZM�/��J��J�	����,ZN�+��}�q��H� �Ιq����Iz�K��Im��z�rO�Lм��4�wU������}0nkl�m�Z�E2�?x���6Q���}��q���ߣ�m�O�f�gAK$�t/��ة;��j%��;�°�i�N8ަ&��խ�����$�7�*�T��l�����h�}+砎=�C-��VZ����+4��6m���fN�T��P6x� 8� �yU�=�/	��[���N?�� f��hh�?\�gϕ���(i�#�G�.��6��@�����ԧHN.��
�I���ۇ�����h�|d�|>�X$� ���>vV�'�6�%c&\	:�:&CiDV�D\*+~�����Ac0��+.��5'����)����^����Lw��h%.tב�h�p<ul�C�B0It�X��H�x1U�t����ޛ�s�b9Ff-7��_aKٲќ}k�Faog��5V��0�{G�V^��+��XZ�\�/I�e����¹Em뼙���
B��|~��O�H�%�
�<M���Ƨ	4k�hi�JWx�4;��j���3�rCq�������^�f���Ӿ���;�|%j��1�p#�z7�ڑ�9nVڲ�=	l�H�D���Q%�oI�'��Oמ6