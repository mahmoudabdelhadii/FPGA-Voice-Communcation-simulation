-- (C) 2001-2016 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
lVTQsct/3AG/3hqIq59N8qO20A1NQDrP1jxdhOpnnoVU+ujCNjcf5XFwYtkUH55rF0r9+9HiCcvQ
ukRqFuemG+EJbI4UKVOJfM5AD9UveRn2pkYy3DcoloeErKJEoQYTsmvhL0jA1rMyVa4EvLZNK/oY
5YuJ/b+/nA94kDhlLFra63ZCt5wzVk5D8evZqAuZ8KUuZQB4dU9UHdWdB2cT60YZC9yylet9b1EH
hzVT0O/RJ7fZ0cQ8tz/IAtdFN6xUHV09PrMc24LSb91q6quIjj5ufxo+feAisC/Ds0sjDdVQ5DDi
wi9cMBy+tENgZbPpWk9m7N98eL1AOPOoog7rXQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 5904)
`protect data_block
ZlK3hWwWf7cR7MKo/qwMxtUm/tlLLzPDYBTTTdfMrUr6PtBibUmuwBGb8wckWzPcJUGGqWRxUvhk
9VKR5FCnHeJ4k0vdU3GPFDLT4QlhsqK0x4+NRUSRNPjX2F3Yfg1AHpcN6RTJo/FrBVwrWUBjHHwl
TRUEm0TcY1GrM+WqPQVYTgUVpkGikQlhOcOPuxeqtXwVUIROJ0Dgw90dRrBhTHGZawyKD0Yl7/AW
YXy38TwLr5Wh6TfoVBqcQmirK8/gmLe+pBfp72aQvwT/h9Mb/QOgi8lAYqx5zDbm1tcajduXeXTu
LJ8KJigONOT4vPWvtPwt3LaGvImneK1lsa+BtMqxGc4G8NvffqVDvVFmokiTdtyqoPNhDzlzdiSN
FeKBiKy7goZN61DqNh4bG/bkwojaHxgHtzTyeX38ZBX8cx6i3OqSIQtbrCSxYInyeaT1nsuPXInR
Be1Vt6kLw8a3ppbb9+buZoj5An/SYXTARflYhhD0yn/rDtaeGJVaPqgdLhZmR5mOdhM7sIxnvu2c
KL685EbsqQx4sMDNYQvUBeVczKHICcdlSqds9Q0RX4vjU3FC1a00orikpcUa3ItCgobtm9KNvz+H
eIddujUQsfStEGpMYNxbGPchWILVdKwMSdcE0rDtC3zZZSkCxhvTjuDFTrQtY7DIbX9b03xjgZAb
XhL9zbAIXoDyLYyGbmiswJ80hV74Q0Tt/7HiW8eyuoYfiBRZwBm67AVl5Q2qaawz+DHSpgCaZxb1
/UKNZcl4RuEhDfi6snEXoFWVHETPpX1q9WzAcrKhOygRv2kxI42QeVd+7N2sRmDuVYtvTa2mhuNV
vz86k/lgrejSrMnuBxXMp+LPVP6T5zmCFO9gYtHn9fpZ2VFxZz0X1Tt/2zAaQS3LM014lwQnGy9z
CMw6uhR9gPb7h601lU/mROEYbTbA9zWBocsS1en+Q0irkHk0EdhE7W3QLr6xNmcGSRaIuyQYg5sd
YjjWYA4Y9guOoEiFHBC2Gs5vlaH5vYPUOTJvOpzoXZ8G7/lVkGc6iJe/dWPLpQnTEJNqGcsUppWJ
woVaVHyscwV22bw4L0h7Ui4NkK35KfC26B4msvG5Np25KItxceTBqs1tvSkfKQxaUp9eufvLyPbW
dsNIBL7E0RwACLB4KVXVZAD1JPIa0X3ZHDs8pfwMUBpxLf1wCt8dm+TPKBR3il5aXFemR3Jg+IyW
UONGUTPyVFZw0nG4PYNOb95pKOuqG6XDjY5QzLGb80G8bjT43S3ch4alibqw+0yvm57lE3H+LfEy
X6PhEYfiCheSZOeClIjzJzg4eTCx8IqEtavb6MG0E6BUDpANC2ndxAJPbzuOYmNUMibHYo1Iq+AL
78CYlR+wwZ9YcI8G3lPLMcPRiBqDlN7Y8wMhMfieuboMdqB/bK4oujFLo0GrEeRNAIYX3/5Vh5/F
h1iMy3aMROpCXcHqfPd4/9N0m927Yp2bwvbfnjby0WCiQTDDZzTAAp0VRPG+Jnyn8naVm2k5bR4k
arZGUlMJeCNJ7GtSrxMNrrxvREv++tEO+CbqTvUPQVC+8HMj1ezPzL6ydKNGscMRh/96JtWAul+E
oOR33YweU1DYnaNssMK2duXhJ6rFaAOT6xx2D0oDx0AjyQWx4U0r5TW4e0xoTOacuoxNA/hcd/tz
igXovKs9iUQkkSjmMDZF2UxI8wxkRbqiOe+n61rQ9pDbLYH3HpXljoO3y6wU+i/hwlSajxToo7d3
ZVroAD0ftvaHZoUwJVDA2TpyejQ4K6hKhKqzoQbuO9aUI2Mjyi3w1p1LhP4UM5fVlURBkAbxczce
OHxmZJZ2RBImJwO2+CXAZPr/V/80BbXgwsKWAhI/l2g8c8lnd0zFPeXkD6rJMiXrGMOsIBisUtmc
TEIjNRajCu+33JK9najMVW9JfrgEw3I95NQOnyFTjROE1mtQdqVoMjx20VPZ5sXCwXgM7X8JLuwF
/dHcLybp10ItjhxPbn5x51wPJxXmvovZh+ZYOV0GNzsAxYzQs89s86Lu21YuSdpe4v8XaKQaYgRC
v1thfJuEx5+L9MVD/UNkyJjRq30S33aHVtbRwFHsYmDZtkpFLccPlxi2TLEVLchMUb1jcoYiHrH8
T/8wYW4QBjUxfeCRexOnVIp7TJjNsLiPR06pZ+0uh95zG8e/yhQWX8ImWVxU/6IWUQDL2Y97ECuP
kor++nPsmZWQrTdy5DwOKny56uvvzf2pgflhHQje7bNpUy6CCfYEn1nj+ZLQ09CDqn2NdoAxEnzH
0iM5i5sXVMRUNjBKXHJlv8Cb007h1eJQa/9KyrLoZgjMozlshQDIG1IDujlocNmhMycaQYwrqOgQ
51UbE8D73VrWGTZHSTfhY26vJ67GWZNYFgiYUqcoBOu0Gkvfa2tdxpELKa9lT2MxAZXr3GF6003m
p5iXSv0aeX26DTpMp7zFHKZcwYn3CI/ScNO3jGyri5XbXLSsl8Uw1sfVIqG0nb9mPmucacBChNEW
YBi5FOO3eqYX+ftfzDsGL7R1iOTX+EUzm9R1kknxAU7hbrqwcJcjHoDSa3R7K+8wcceCFbMmuFYe
vU2tQlEkSYI1HzcaeQF0AGkcCmru00VlxfClk3RZfBDb5m/mK2GQpVS6yTFQjuHmg0MXNtmnkrQv
DPRBrrdSWnazK1ugyf7Hi/GANcqIESeajCe3KBmzz+wv2PzBy+Zf5N3XCMyP/fhKfb9QhRke3rSc
jcc7PGGB7w7KP0V+KccMqk28vCMheCn9FIkGViuD5K8mlZYk3EjLGOy89rTcKS3hQ2A4YRGdjyG8
EZtroNd8bzScPlrn+08eoQiUq/q6xcaXo2ZAIO3heSRtaXgeyBqgKyglNKnS9ij0ktmnYq93RutH
Oe7tiyri5fNZpwyeHkdaBmE/rHBaW/8DgsSwCKrAwoUW17KFZl4dJ945Px3GChtkbL8xlADrhPPO
nXc7U/cXj6g3HD2Lt9xvCu3oY1t9562zeGRWufBTLyB957o5vaQZqEevo+WnsfuOa6cXuwShXjsL
uk883w3eOlslfmjOP8tgZqYqN5q5ouCOMH0sEUsSjE2ZJGateJ7smIY33nLJGig4F8w67HDNV0aL
cR2JXyHNpfgmBiTrlWliQMj+HXI0t0TuZM5RWM7YYavuFMuda4YpuhC9VfX4uQtQYSVSnv9yz+dj
9827TufzL/K9Hz6WixIMcC8hp2eFBKObEHGo7RcwHp+EQoI2a8PlpWcRSegLH1w/gzhtAObpnwn6
iKdltxJEwpfi7sU7GaSj2rhePLY7if4cay3y8QGLeryuZu8W68s9vWv3k2ofNG4LoSa76jEVEqRv
dKE18z4J/BNL4TWOm0nyKHjcmxML7DFguwhhCq3mb3ZEJRYXG+o6gCUi4KCUrA0VJdbx8lTqmUtc
TutSs2p2O+ni+GozL2HxYhkgJ/CdO4zIck988VEt8C8QwcE9Cl6EPJu/cgUoH8jW2OLTjPIZdr7t
mWM6uF/EvTej/F8nd+GwHip0reUoN6I9m8wWZkcjU+xKdMO2dmDdiyhYr5dcveEDxtDNLn5y18iF
7G5AbwC/GFVc4nnizlDdb9vuU3GMnhm8TqRFagiUAmnYBD9KmEP1/s5U0qxkBy0eLlWwMzGFlRzt
Q9H+8qpJuHSr628DaM/4DOmXbkwCayc+GcSBzXVGM6MCfBPGHLVcMKc+5mppyw/uNCLm8ILMtC25
cyrStu6pc12a+qkDyWbhPrHdfwRmHf43QR7sZRSOXRNG+Xqj0lIrve+ZysbJBKAofsc1AukwElyJ
Nl3p0Nh3DWPPns/UbBzl4nL1+0Oy1FkiKOpTMEiMjbvlduyivmxLlh7GZeJrrFjRMu+f8GlRugb5
0GItzEohJ/vOI3MF8tNkw4PRGKk1RamDC/chyHkiwpDXTB230DJZdHrcsE/TnGtzQw8h8BtebKXQ
dvvFGxWog00+203yDyVoRXO8ApDSTEpWCmyLxBulzzRB8sdQmenjduYlPgNm5/yOFPPGaYxzqWHu
lKMwpjHTf30+iqoYK+ltw7D9srXZ+QpgB1L95VV/frOg0irKPy6SPSmws912U1yQuO+yYVUesp6p
vh8jZ5YTUfuIGefmkADT+2L3ZvU5ab+0YTIFFnJA+tuuyimuWJuOJd6zZlf6z5dGh7yNy9PT5j76
JfauuAtZ03UD0G62VxmWxIvqP8KYWA0x/aYYTniL7Zl6nHe81mAnyeO0aMSPpLahhQQE8Bok0sRB
8fHNKt71xyPQfSwjN9+gCEEhvglalx1H/xhZaf4TFbOTzqb1FwTVxnFq7FYWktuYakKTZGOo5UaM
XVNDsTdI02FUnxYGaGVmuoWy29budbirGH8djberewDhzAxZzv6gZTGKRTHc2Wk55kJ1zEZ8vTSY
YQm7IsCIJNkeTpaYo2j3+DmNhc0cwgTVK48Uc2Of29Vk9toTOXvYPnwgkjHUcmxhVyKfTbqxQinZ
0reXU0dEvLUFVnVmsUMaRRilo21dZcGYwjn3Yxux7sVIJPGuLKvysBfWMt3QjpfujQGtmq6JkIlF
vwL8IXtkHFMzbHpe3ouUloy7ZNNB38F0s33WXvRGq1yLmoQKuNtx0tq8UJB3eqntGMGuCbg824PZ
nksb5S5VYZquJYjuAn880hPolcQR0bveiBeYoQgHKesbJFuldPK9tlClTk6gC6QFsz/oSe2PM5jq
UnixxOlkLV8kuHxhb3Igi9uYf07D1u6AmpYUEhPehYX7nyCyPwJsK1eOFmBTN2mdpYsOUNx7FjP+
WX3VPsBWFQXYhUQtdgIYlFjck2v3NFPBnvGEA3363RjQV2JX6k+hcvZwYNKLAKw7UIhLwxBzpPio
cgSvfVXKs+iyJ27hKSO9NiaqSqTg4YA1tMbkg4ukVgGrdEminM9S2s+BhhzAzHisC2EXLUpdLWt+
YwWDa0E6r9bWlT0hnELmDuRWOL30HyR8FAt0Hk6joOaZsAfrgciiagshoXQIcbRcL0i9cbvAMJIn
7uulUek6Z7M2SYMM6oWEYgtPa/oj0g0PmS0OcI/DrAvHOR5HYtdbDkrXH88vQq82D9TW2MgoaeXa
4En+Pth89TxWjSD2/+DFcpN999Ng+KoGr5l6/K+qQirJwuLCff0X4OXIGvGiAPSgRz8oFqpXlkKd
6hRq327rVBPBpPcqegXOO5PZanYOOcN2CwxfN82a/5xxr/ea1nN6O+D+va4KtngJXGLBeCiDrKOD
x/jeCfo8QoomodJG7cO1U/O51GiSZo27t9SJ90ngX8vt0nlY6gQMkRqIHMRgslWbZKyan0dgB8nM
MXDB7S7Y4Op2r6J6aNoSQKsHMybXnEHEiF/9Djj2jGkOgFwqFDEIECtPYI9bKZ+JSDYpN27hn/es
uWrQ7hqLbrtWFxFnnrK9f0v1YCHtYyfWHIj0o64CefaRvT9HjXRUeL2m6x+TujBVm0zFK0fGUnFG
FhVxNRRNM0UayIhXVFGZtGzQnQSLndBLbyrF2ZOBP3PWiy1D2L5BTvBkPP7aW8pF2O+D4dSgdcsF
zCYkl6/jz5yFDpZ38ynirAJOGV1QRKvmaox7iYkr5nxujwsPyDIP8HgZumHau6iIcyMtFOmOBzk9
N1cXKrUs+EaToXiidVse6vp8U1GJs1mle92ZuFLwCwcOuVKcMoNZV/ehyF8X5Yeabq1AbY7eRY4n
ThNDrdWhLU+b6uIq2b6UFJnwgK39vKqZ9elFsSnuQE5N40M22HQpTG3AdsFik+uiP/UjqSBNSzKX
7z8LWfZu00TTfLuHhqiCrbcCssRBIu1+RQNewwdQvrUexfrRRlnEKJUfKXdP8Tto8WCsbOcCQR37
BrDKVaoAZogBmuMXVswe/dxxDuXIfaOtSPRbUv/pDyIiKoNdlqnvgKy6WeVz1ww6j35W5ZrgPtCX
HZpyuOVId5XkipLSncvNpW0tpWheF4tW9I+4AAQoVQdx4oqxpeT6BkELqbYMjfUUBSgs4FfyW1bU
0PF4l5nxuxyWEwz3tSQKbiDJRBAb/50jV5hbjbDVjwscDs63xZFy0hMo/SNixXRlTB89hVZfJ65s
abF+THbL5mERo1s7E6WcNIF8h8MOWJ5svMPpcI/jx0Y7Y+Ar2rvWQ5cwpnY972yanmM+J9n7oD/4
3vi63OEmC9wOf8YWbJ1C7IVCAmKCocVWpHLB0g5gSG9YLKnCJw2J3eB+ejOx1qWDtEKlOw5BaerU
O+gjUmDpBVhHYtCaKxjSR8dWmcHrmzRTFO+e68hyE6p5dIh1Kr1g/Eb/Iw+wHOUblCWihOSoudcA
7OFdaxEYhXu0A+PzDOpg5FC0rZbMR/kSNcEBqXWmSSHVZaSXY2sWvIbwS/EOpkFjuqr6TkAf3xlj
uRgZ0U/UXvCY16YFJ2qR8NKiItIRdAE7dKRxawgKp8oxksisRd763A0I0DprKm6SfH/L9xjaTi1T
Ci2wEWHpF7ZCfA1kGOjM/UBf5cvo0uvUtjJwgrr5yQdoLAe59ty5xgiKdt6FIrUx4xMMQW7f6YaP
qxVksxqW7te6LO9q5SRXdzwqHmrifnSsPPqrWetGWrHvFnGjpwcH+E2xy0f1wCl+QkAp3sdY1VRo
mkwS4BlZZ6V1yFLn5EQNR1TbT2YRwU/LIRjZG8L0/ZOcLQzbmI0PrOyfSj62VP/e4kutIYppIxD8
jZ3g/fnEktg0i/3twQkxHnds+wCH5J3Fz7VHgYSIRHxSHwt4+dR2DeosMpFlW1NIDAQbcln8ddA3
ASqBpA2fQHeYxcMTW9GI95LpyfF5gBbE6Ll4As75IGvQiSv2VNYz2Dj+p3PoCBAfn73vy7xUG5i5
oSGY/0+DpT5sODG/RuW0BuptTcMXErV2J2f12IkndI8IweQFtsgcm/MSUq3tcrfLtXgo7Ed+I3gw
6GDAarEl8SMB8E/kqFDEupq4xoNuNPIXcxGtFcSznhW6Y4FYKQRrJSPD0eM1Hq0+zNT0v+sD6U95
7/7h1ZcUGCa01q/rbi9P2cI+x4YhKaQRG9NqynDsAcYqgtAbUz6J2qNoTx8/00O7GXeed8tAokgl
4PNQa6Gc3kpnpkz2ahow06Q7OfZtwllYI9UvLsbP5HQBkUk5N5/11wD3lxJdzEEpa6oeAZPVZeBe
GQk35+lgNK2W64qmWkAIY1Ade7OzJHMiz8iXmfuMu39PVxhb4zhnk/WBmWqj8ufAzaRE10AB5uhc
uzDf16j+O+2Z11jihyfyPR+0oMkbxudaYGnigP4CKteZiD8wVUSb8NR6Pu1Q20sN8kURBddKhv1R
CPydbUy85VuhhN9kg9xWdvZpYg3zv0W1QMExhA58esHcaewvrk87oFXfNgr8p3twaTuklginVqLt
+7igfaxpFZm2ODYRM0AXLwEmT2OP85/a0kr7mj7/IlXN6wx82mexeCd/qInKtk8I7LJQ3SY7en8X
6j/rj2/0dPdjBYvJgVWtda1EHO2ORXEgfUWkLzUGlsCDSZ33SOx8AusqPQX2+uDM/OpH6lpssrUI
A4o0k+av+utCOqgiEekG8IG2CoIZ2yrtpPyEz9+yvhmi6t9XDQ/TUrMMjM5tQA4sxf0IQppWtir1
aEaByoQ2oJV6fr7U8k9de8BzH4SnGhRwOTJFp/vNqlWqEIssuiiNczAwbEER5AP7Qn028UZu6sVH
FTYi5mH0G1SGXaHdWHh5HOj65pqv5jvYakSTf2F9fzxxWC0pVeFVclqkQS59hZlo9cj45rUWIF34
8jS0Ym9E3N5Ho5mODlXRHZgoV/5koySQx+kuXJXZRK+ZJgej8dqtXZIzh/8JMSGLEszZGR6JRps5
Q7xYEsHyLZmbbFrEX6Wp1F1dsArJmdRJ0aHCmnzTIdRI
`protect end_protected
